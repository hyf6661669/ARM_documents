VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;

SITE TSM90NMADSITE
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE 0.280 BY 2.520 ;
END TSM90NMADSITE

MACRO ACCSHCINX2AD
    CLASS CORE ;
    FOREIGN ACCSHCINX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.945 1.425 7.065 1.820 ;
        RECT  6.730 1.425 6.945 1.655 ;
        RECT  6.560 0.870 6.730 1.655 ;
        RECT  6.305 1.425 6.560 1.655 ;
        RECT  6.185 1.425 6.305 1.835 ;
        END
        AntennaDiffArea 0.378 ;
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.145 1.780 8.265 2.040 ;
        RECT  8.090 1.285 8.145 2.115 ;
        RECT  8.025 0.720 8.090 2.115 ;
        RECT  7.885 0.720 8.025 1.420 ;
        RECT  7.545 1.995 8.025 2.115 ;
        RECT  7.425 1.780 7.545 2.115 ;
        END
        AntennaDiffArea 0.417 ;
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.030 1.010 9.170 1.655 ;
        END
        AntennaGateArea 0.147 ;
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.650 0.905 8.890 1.375 ;
        END
        AntennaGateArea 0.147 ;
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 1.115 3.595 1.375 ;
        RECT  2.910 1.195 3.430 1.315 ;
        RECT  2.740 1.195 2.910 1.365 ;
        END
        AntennaGateArea 0.403 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 1.125 0.490 1.375 ;
        END
        AntennaGateArea 0.147 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.075 -0.210 9.520 0.210 ;
        RECT  8.865 -0.210 9.075 0.460 ;
        RECT  5.115 -0.210 8.865 0.210 ;
        RECT  4.855 -0.210 5.115 0.370 ;
        RECT  1.055 -0.210 4.855 0.210 ;
        RECT  0.885 -0.210 1.055 0.315 ;
        RECT  0.635 -0.210 0.885 0.210 ;
        RECT  0.465 -0.210 0.635 0.735 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.025 2.310 9.520 2.730 ;
        RECT  8.905 1.800 9.025 2.730 ;
        RECT  5.115 2.310 8.905 2.730 ;
        RECT  4.855 2.285 5.115 2.730 ;
        RECT  1.310 2.310 4.855 2.730 ;
        RECT  1.050 2.220 1.310 2.730 ;
        RECT  0.255 2.310 1.050 2.730 ;
        RECT  0.085 1.770 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.520 2.520 ;
        LAYER M1 ;
        RECT  9.315 0.415 9.435 2.155 ;
        RECT  9.265 0.415 9.315 0.845 ;
        RECT  9.290 1.635 9.315 2.155 ;
        RECT  8.735 0.605 9.265 0.725 ;
        RECT  8.615 0.390 8.735 0.725 ;
        RECT  8.385 1.525 8.625 2.090 ;
        RECT  6.200 0.390 8.615 0.510 ;
        RECT  8.385 0.700 8.485 0.820 ;
        RECT  8.265 0.700 8.385 1.660 ;
        RECT  8.225 0.700 8.265 0.820 ;
        RECT  7.785 1.540 7.905 1.870 ;
        RECT  7.545 1.540 7.785 1.660 ;
        RECT  7.545 0.630 7.730 0.750 ;
        RECT  7.425 0.630 7.545 1.660 ;
        RECT  6.440 0.630 7.425 0.750 ;
        RECT  7.185 0.895 7.305 2.140 ;
        RECT  6.880 0.895 7.185 1.015 ;
        RECT  6.755 2.020 7.185 2.140 ;
        RECT  6.495 1.800 6.755 2.140 ;
        RECT  1.625 2.020 6.495 2.140 ;
        RECT  6.320 0.630 6.440 1.200 ;
        RECT  5.950 1.080 6.320 1.200 ;
        RECT  6.080 0.390 6.200 0.960 ;
        RECT  5.805 0.815 6.080 0.960 ;
        RECT  5.825 1.375 5.945 1.900 ;
        RECT  5.805 1.375 5.825 1.495 ;
        RECT  5.675 0.815 5.805 1.495 ;
        RECT  5.575 0.415 5.745 0.610 ;
        RECT  5.565 1.640 5.685 1.900 ;
        RECT  4.655 0.490 5.575 0.610 ;
        RECT  2.000 1.780 5.565 1.900 ;
        RECT  5.425 1.100 5.530 1.360 ;
        RECT  5.425 0.805 5.450 0.975 ;
        RECT  5.305 0.805 5.425 1.660 ;
        RECT  5.280 0.805 5.305 0.975 ;
        RECT  5.000 1.145 5.170 1.315 ;
        RECT  4.690 1.145 5.000 1.265 ;
        RECT  4.685 1.145 4.690 1.615 ;
        RECT  4.520 0.745 4.685 1.615 ;
        RECT  4.530 0.380 4.655 0.610 ;
        RECT  4.095 0.380 4.530 0.500 ;
        RECT  4.515 0.745 4.520 1.470 ;
        RECT  4.255 0.745 4.515 0.915 ;
        RECT  4.280 1.540 4.370 1.660 ;
        RECT  4.160 1.050 4.280 1.660 ;
        RECT  4.095 1.050 4.160 1.180 ;
        RECT  3.325 1.540 4.160 1.660 ;
        RECT  3.975 0.380 4.095 1.180 ;
        RECT  3.035 0.380 3.975 0.500 ;
        RECT  3.835 1.300 3.975 1.420 ;
        RECT  3.715 0.620 3.835 1.420 ;
        RECT  2.885 0.620 3.715 0.740 ;
        RECT  2.620 1.540 3.205 1.660 ;
        RECT  2.760 0.385 2.885 0.740 ;
        RECT  2.620 0.865 2.800 0.985 ;
        RECT  1.300 0.385 2.760 0.505 ;
        RECT  2.500 0.625 2.620 1.660 ;
        RECT  1.540 0.625 2.500 0.745 ;
        RECT  2.200 1.540 2.500 1.660 ;
        RECT  2.000 0.865 2.380 0.985 ;
        RECT  1.880 0.865 2.000 1.900 ;
        RECT  1.430 1.470 1.690 1.850 ;
        RECT  1.505 1.980 1.625 2.140 ;
        RECT  1.420 0.625 1.540 1.290 ;
        RECT  1.060 1.980 1.505 2.100 ;
        RECT  1.300 1.470 1.430 1.620 ;
        RECT  1.180 0.385 1.300 1.620 ;
        RECT  0.925 0.640 1.060 2.100 ;
        RECT  0.800 0.640 0.925 0.760 ;
        RECT  0.715 1.930 0.925 2.100 ;
        RECT  0.645 0.880 0.805 1.755 ;
        RECT  0.255 0.880 0.645 1.000 ;
        RECT  0.470 1.495 0.645 1.755 ;
        RECT  0.085 0.475 0.255 1.000 ;
    END
END ACCSHCINX2AD
MACRO ACCSHCINX4AD
    CLASS CORE ;
    FOREIGN ACCSHCINX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.915 1.275 7.080 1.820 ;
        RECT  6.775 1.275 6.915 1.430 ;
        RECT  6.515 0.880 6.775 1.430 ;
        RECT  6.370 1.275 6.515 1.430 ;
        RECT  6.200 1.275 6.370 1.835 ;
        END
        AntennaDiffArea 0.361 ;
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.160 1.750 8.280 2.010 ;
        RECT  8.040 0.680 8.160 2.140 ;
        RECT  7.910 0.680 8.040 1.235 ;
        RECT  7.560 2.020 8.040 2.140 ;
        RECT  7.440 1.780 7.560 2.140 ;
        END
        AntennaDiffArea 0.355 ;
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.030 1.015 9.170 1.515 ;
        END
        AntennaGateArea 0.1483 ;
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.670 1.030 8.890 1.375 ;
        END
        AntennaGateArea 0.1482 ;
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 1.115 3.595 1.375 ;
        RECT  2.910 1.195 3.430 1.315 ;
        RECT  2.740 1.195 2.910 1.365 ;
        END
        AntennaGateArea 0.3859 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 1.125 0.490 1.375 ;
        END
        AntennaGateArea 0.148 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.040 -0.210 9.520 0.210 ;
        RECT  8.780 -0.210 9.040 0.390 ;
        RECT  5.090 -0.210 8.780 0.210 ;
        RECT  4.830 -0.210 5.090 0.370 ;
        RECT  1.055 -0.210 4.830 0.210 ;
        RECT  0.885 -0.210 1.055 0.315 ;
        RECT  0.635 -0.210 0.885 0.210 ;
        RECT  0.465 -0.210 0.635 0.735 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.025 2.310 9.520 2.730 ;
        RECT  8.855 1.845 9.025 2.730 ;
        RECT  5.090 2.310 8.855 2.730 ;
        RECT  4.830 2.285 5.090 2.730 ;
        RECT  1.310 2.310 4.830 2.730 ;
        RECT  1.050 2.220 1.310 2.730 ;
        RECT  0.255 2.310 1.050 2.730 ;
        RECT  0.085 1.770 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.520 2.520 ;
        LAYER M1 ;
        RECT  9.290 0.380 9.410 2.180 ;
        RECT  9.240 0.380 9.290 0.900 ;
        RECT  9.215 1.750 9.290 2.180 ;
        RECT  8.415 0.510 9.240 0.630 ;
        RECT  8.490 1.495 8.640 2.140 ;
        RECT  8.490 0.750 8.630 0.870 ;
        RECT  8.400 0.750 8.490 2.140 ;
        RECT  8.295 0.390 8.415 0.630 ;
        RECT  8.370 0.750 8.400 1.655 ;
        RECT  6.155 0.390 8.295 0.510 ;
        RECT  7.800 1.500 7.920 1.900 ;
        RECT  7.650 1.500 7.800 1.620 ;
        RECT  7.650 0.710 7.760 0.970 ;
        RECT  7.530 0.630 7.650 1.620 ;
        RECT  6.395 0.630 7.530 0.750 ;
        RECT  7.200 0.880 7.320 2.060 ;
        RECT  6.895 0.880 7.200 1.000 ;
        RECT  6.700 1.940 7.200 2.060 ;
        RECT  6.580 1.670 6.700 2.140 ;
        RECT  1.625 2.020 6.580 2.140 ;
        RECT  6.275 0.630 6.395 1.130 ;
        RECT  5.915 1.010 6.275 1.130 ;
        RECT  6.035 0.390 6.155 0.850 ;
        RECT  5.795 0.730 6.035 0.850 ;
        RECT  5.840 1.375 5.960 1.900 ;
        RECT  5.745 0.415 5.915 0.610 ;
        RECT  5.795 1.375 5.840 1.495 ;
        RECT  5.675 0.730 5.795 1.495 ;
        RECT  4.630 0.490 5.745 0.610 ;
        RECT  5.560 1.640 5.680 1.900 ;
        RECT  2.000 1.780 5.560 1.900 ;
        RECT  5.400 1.100 5.555 1.360 ;
        RECT  5.400 0.805 5.425 0.975 ;
        RECT  5.280 0.805 5.400 1.660 ;
        RECT  5.255 0.805 5.280 0.975 ;
        RECT  4.975 1.145 5.145 1.315 ;
        RECT  4.665 1.145 4.975 1.265 ;
        RECT  4.660 1.145 4.665 1.615 ;
        RECT  4.490 0.745 4.660 1.615 ;
        RECT  4.505 0.380 4.630 0.610 ;
        RECT  4.095 0.380 4.505 0.500 ;
        RECT  4.215 0.745 4.490 0.915 ;
        RECT  4.280 1.540 4.370 1.660 ;
        RECT  4.160 1.050 4.280 1.660 ;
        RECT  4.095 1.050 4.160 1.180 ;
        RECT  3.325 1.540 4.160 1.660 ;
        RECT  3.975 0.380 4.095 1.180 ;
        RECT  3.035 0.380 3.975 0.500 ;
        RECT  3.835 1.300 3.975 1.420 ;
        RECT  3.715 0.620 3.835 1.420 ;
        RECT  2.885 0.620 3.715 0.740 ;
        RECT  2.620 1.540 3.205 1.660 ;
        RECT  2.760 0.385 2.885 0.740 ;
        RECT  2.620 0.865 2.800 0.985 ;
        RECT  1.300 0.385 2.760 0.505 ;
        RECT  2.500 0.625 2.620 1.660 ;
        RECT  1.540 0.625 2.500 0.745 ;
        RECT  2.200 1.540 2.500 1.660 ;
        RECT  2.000 0.865 2.380 0.985 ;
        RECT  1.880 0.865 2.000 1.900 ;
        RECT  1.430 1.470 1.690 1.850 ;
        RECT  1.505 1.980 1.625 2.140 ;
        RECT  1.420 0.625 1.540 1.290 ;
        RECT  1.060 1.980 1.505 2.100 ;
        RECT  1.300 1.470 1.430 1.620 ;
        RECT  1.180 0.385 1.300 1.620 ;
        RECT  0.925 0.640 1.060 2.100 ;
        RECT  0.800 0.640 0.925 0.760 ;
        RECT  0.715 1.930 0.925 2.100 ;
        RECT  0.685 0.880 0.805 1.755 ;
        RECT  0.255 0.880 0.685 1.000 ;
        RECT  0.470 1.495 0.685 1.755 ;
        RECT  0.085 0.475 0.255 1.000 ;
    END
END ACCSHCINX4AD
MACRO ACCSHCONX2AD
    CLASS CORE ;
    FOREIGN ACCSHCONX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.300 0.620 6.420 1.220 ;
        RECT  5.530 0.620 6.300 0.740 ;
        RECT  6.125 1.100 6.300 1.220 ;
        RECT  6.005 1.100 6.125 1.785 ;
        RECT  5.510 0.620 5.530 1.095 ;
        RECT  5.390 0.620 5.510 1.650 ;
        RECT  5.215 1.530 5.390 1.650 ;
        END
        AntennaDiffArea 0.479 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.190 1.615 7.360 1.900 ;
        RECT  7.060 0.665 7.230 1.265 ;
        RECT  6.930 1.615 7.190 1.735 ;
        RECT  6.930 1.145 7.060 1.265 ;
        RECT  6.790 1.145 6.930 1.735 ;
        RECT  6.615 1.615 6.790 1.735 ;
        RECT  6.495 1.615 6.615 1.895 ;
        END
        AntennaDiffArea 0.425 ;
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.175 0.995 8.330 1.425 ;
        END
        AntennaGateArea 0.162 ;
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.860 1.045 8.050 1.415 ;
        RECT  7.680 1.045 7.860 1.215 ;
        END
        AntennaGateArea 0.162 ;
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.915 0.910 3.345 1.235 ;
        RECT  2.825 0.910 2.915 1.095 ;
        END
        AntennaGateArea 0.4626 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.045 0.320 1.215 ;
        RECT  0.070 1.045 0.210 1.655 ;
        END
        AntennaGateArea 0.3233 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.065 -0.210 8.680 0.210 ;
        RECT  7.805 -0.210 8.065 0.390 ;
        RECT  4.680 -0.210 7.805 0.210 ;
        RECT  4.510 -0.210 4.680 0.705 ;
        RECT  3.655 -0.210 4.510 0.210 ;
        RECT  3.485 -0.210 3.655 0.550 ;
        RECT  1.330 -0.210 3.485 0.210 ;
        RECT  1.070 -0.210 1.330 0.390 ;
        RECT  0.265 -0.210 1.070 0.210 ;
        RECT  0.100 -0.210 0.265 0.875 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.080 2.310 8.680 2.730 ;
        RECT  7.910 1.610 8.080 2.730 ;
        RECT  4.340 2.310 7.910 2.730 ;
        RECT  4.080 2.210 4.340 2.730 ;
        RECT  3.505 2.310 4.080 2.730 ;
        RECT  3.335 2.265 3.505 2.730 ;
        RECT  1.310 2.310 3.335 2.730 ;
        RECT  1.050 2.170 1.310 2.730 ;
        RECT  0.260 2.310 1.050 2.730 ;
        RECT  0.100 1.800 0.260 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.680 2.520 ;
        LAYER M1 ;
        RECT  8.465 0.520 8.570 1.675 ;
        RECT  8.450 0.520 8.465 2.065 ;
        RECT  8.280 0.400 8.450 0.830 ;
        RECT  8.295 1.545 8.450 2.065 ;
        RECT  7.635 0.520 8.280 0.640 ;
        RECT  7.550 1.375 7.720 1.990 ;
        RECT  7.480 0.760 7.655 0.880 ;
        RECT  7.515 0.380 7.635 0.640 ;
        RECT  7.480 1.375 7.550 1.495 ;
        RECT  5.270 0.380 7.515 0.500 ;
        RECT  7.360 0.760 7.480 1.495 ;
        RECT  6.905 1.855 7.045 1.975 ;
        RECT  6.785 1.855 6.905 2.140 ;
        RECT  6.660 0.715 6.870 0.995 ;
        RECT  6.375 2.020 6.785 2.140 ;
        RECT  6.540 0.715 6.660 1.495 ;
        RECT  6.375 1.360 6.540 1.495 ;
        RECT  6.255 1.360 6.375 2.140 ;
        RECT  4.575 2.015 6.255 2.140 ;
        RECT  5.850 0.860 6.110 0.980 ;
        RECT  5.730 0.860 5.850 1.895 ;
        RECT  5.645 1.550 5.730 1.895 ;
        RECT  4.790 1.775 5.645 1.895 ;
        RECT  5.150 0.330 5.270 1.345 ;
        RECT  5.080 1.225 5.150 1.345 ;
        RECT  4.960 1.225 5.080 1.655 ;
        RECT  4.900 1.485 4.960 1.655 ;
        RECT  4.815 0.520 4.935 1.040 ;
        RECT  4.705 0.825 4.815 1.040 ;
        RECT  4.670 1.730 4.790 1.895 ;
        RECT  4.585 0.825 4.705 1.610 ;
        RECT  4.375 1.730 4.670 1.850 ;
        RECT  4.295 0.825 4.585 0.945 ;
        RECT  4.475 1.970 4.575 2.140 ;
        RECT  3.555 1.970 4.475 2.090 ;
        RECT  4.255 1.090 4.375 1.850 ;
        RECT  4.175 0.675 4.295 0.945 ;
        RECT  3.895 1.090 4.255 1.210 ;
        RECT  4.015 1.330 4.135 1.850 ;
        RECT  3.895 0.375 4.015 0.545 ;
        RECT  3.270 1.730 4.015 1.850 ;
        RECT  3.775 0.375 3.895 1.610 ;
        RECT  3.715 1.440 3.775 1.610 ;
        RECT  3.465 0.670 3.585 1.610 ;
        RECT  3.435 1.970 3.555 2.140 ;
        RECT  3.295 0.670 3.465 0.790 ;
        RECT  3.030 1.490 3.465 1.610 ;
        RECT  1.615 2.020 3.435 2.140 ;
        RECT  3.125 0.355 3.295 0.790 ;
        RECT  3.150 1.730 3.270 1.900 ;
        RECT  1.930 1.780 3.150 1.900 ;
        RECT  2.800 0.670 3.125 0.790 ;
        RECT  2.910 1.490 3.030 1.660 ;
        RECT  2.170 1.540 2.910 1.660 ;
        RECT  2.580 0.380 2.870 0.525 ;
        RECT  2.580 1.300 2.810 1.420 ;
        RECT  2.460 0.380 2.580 1.420 ;
        RECT  1.570 0.380 2.460 0.500 ;
        RECT  1.930 0.625 2.295 0.795 ;
        RECT  2.050 1.330 2.170 1.660 ;
        RECT  1.810 0.625 1.930 1.900 ;
        RECT  1.650 0.760 1.690 0.880 ;
        RECT  1.530 0.760 1.650 1.810 ;
        RECT  1.495 1.930 1.615 2.140 ;
        RECT  1.450 0.380 1.570 0.640 ;
        RECT  1.430 0.760 1.530 0.880 ;
        RECT  1.475 1.380 1.530 1.810 ;
        RECT  0.615 1.930 1.495 2.050 ;
        RECT  0.915 0.520 1.450 0.640 ;
        RECT  1.290 1.000 1.410 1.260 ;
        RECT  0.885 1.025 1.290 1.195 ;
        RECT  0.885 0.375 0.915 0.640 ;
        RECT  0.765 0.375 0.885 1.670 ;
        RECT  0.715 1.500 0.765 1.670 ;
        RECT  0.565 0.720 0.615 0.890 ;
        RECT  0.565 1.930 0.615 2.100 ;
        RECT  0.445 0.720 0.565 2.100 ;
    END
END ACCSHCONX2AD
MACRO ACCSHCONX4AD
    CLASS CORE ;
    FOREIGN ACCSHCONX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.700 0.620 6.850 0.740 ;
        RECT  6.580 0.620 6.700 1.220 ;
        RECT  5.820 0.620 6.580 0.740 ;
        RECT  6.570 1.100 6.580 1.220 ;
        RECT  6.450 1.100 6.570 1.785 ;
        RECT  5.820 1.540 5.920 1.660 ;
        RECT  5.670 0.620 5.820 1.660 ;
        RECT  5.160 1.540 5.670 1.660 ;
        RECT  5.020 0.450 5.160 1.660 ;
        RECT  4.900 1.480 5.020 1.600 ;
        END
        AntennaDiffArea 0.78 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.450 1.660 8.590 1.780 ;
        RECT  8.320 1.660 8.450 2.140 ;
        RECT  8.195 0.750 8.350 0.870 ;
        RECT  7.805 2.010 8.320 2.140 ;
        RECT  8.075 0.620 8.195 0.870 ;
        RECT  7.525 0.620 8.075 0.740 ;
        RECT  7.675 1.605 7.805 2.140 ;
        RECT  7.525 1.605 7.675 1.735 ;
        RECT  7.350 0.620 7.525 1.735 ;
        RECT  7.080 1.605 7.350 1.735 ;
        RECT  6.960 1.605 7.080 1.895 ;
        END
        AntennaDiffArea 0.735 ;
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.450 1.020 9.675 1.375 ;
        RECT  9.310 0.865 9.450 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.610 1.085 8.925 1.255 ;
        RECT  8.470 0.865 8.610 1.255 ;
        END
        AntennaGateArea 0.324 ;
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.130 3.390 1.375 ;
        RECT  3.070 1.130 3.150 1.250 ;
        END
        AntennaGateArea 0.4644 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 1.045 0.395 1.215 ;
        RECT  0.070 1.045 0.240 1.655 ;
        END
        AntennaGateArea 0.3233 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.205 -0.210 10.360 0.210 ;
        RECT  10.050 -0.210 10.205 0.885 ;
        RECT  9.535 -0.210 10.050 0.210 ;
        RECT  9.275 -0.210 9.535 0.390 ;
        RECT  8.675 -0.210 9.275 0.210 ;
        RECT  8.555 -0.210 8.675 0.380 ;
        RECT  4.695 -0.210 8.555 0.210 ;
        RECT  4.525 -0.210 4.695 0.520 ;
        RECT  3.675 -0.210 4.525 0.210 ;
        RECT  3.530 -0.210 3.675 0.645 ;
        RECT  1.360 -0.210 3.530 0.210 ;
        RECT  1.100 -0.210 1.360 0.390 ;
        RECT  0.255 -0.210 1.100 0.210 ;
        RECT  0.085 -0.210 0.255 0.840 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.255 2.310 10.360 2.730 ;
        RECT  10.085 1.555 10.255 2.730 ;
        RECT  9.535 2.310 10.085 2.730 ;
        RECT  9.365 1.565 9.535 2.730 ;
        RECT  8.815 2.310 9.365 2.730 ;
        RECT  8.645 1.980 8.815 2.730 ;
        RECT  4.390 2.310 8.645 2.730 ;
        RECT  4.130 2.210 4.390 2.730 ;
        RECT  3.600 2.310 4.130 2.730 ;
        RECT  3.340 2.260 3.600 2.730 ;
        RECT  1.380 2.310 3.340 2.730 ;
        RECT  1.120 2.190 1.380 2.730 ;
        RECT  0.255 2.310 1.120 2.730 ;
        RECT  0.085 1.845 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.360 2.520 ;
        LAYER M1 ;
        RECT  9.805 0.405 9.930 1.995 ;
        RECT  9.680 0.405 9.805 0.835 ;
        RECT  9.725 1.565 9.805 1.995 ;
        RECT  8.435 0.510 9.680 0.630 ;
        RECT  9.045 0.760 9.175 1.995 ;
        RECT  8.915 0.760 9.045 0.880 ;
        RECT  9.005 1.375 9.045 1.995 ;
        RECT  8.185 1.375 9.005 1.495 ;
        RECT  8.315 0.380 8.435 0.630 ;
        RECT  5.550 0.380 8.315 0.500 ;
        RECT  8.015 1.335 8.185 1.890 ;
        RECT  7.950 1.335 8.015 1.455 ;
        RECT  7.830 0.860 7.950 1.455 ;
        RECT  7.690 0.860 7.830 0.980 ;
        RECT  7.370 1.855 7.510 1.975 ;
        RECT  7.250 1.855 7.370 2.140 ;
        RECT  6.840 2.020 7.250 2.140 ;
        RECT  6.995 0.715 7.165 1.460 ;
        RECT  6.840 1.340 6.995 1.460 ;
        RECT  6.720 1.340 6.840 2.140 ;
        RECT  4.630 2.020 6.720 2.140 ;
        RECT  6.210 0.860 6.460 0.980 ;
        RECT  6.090 0.860 6.210 1.900 ;
        RECT  4.875 1.780 6.090 1.900 ;
        RECT  5.430 0.380 5.550 1.420 ;
        RECT  5.280 1.300 5.430 1.420 ;
        RECT  4.860 0.755 4.885 0.935 ;
        RECT  4.755 1.725 4.875 1.900 ;
        RECT  4.750 0.720 4.860 0.980 ;
        RECT  4.480 1.725 4.755 1.845 ;
        RECT  4.740 0.720 4.750 1.600 ;
        RECT  4.715 0.755 4.740 1.600 ;
        RECT  4.630 0.815 4.715 1.600 ;
        RECT  4.310 0.815 4.630 0.935 ;
        RECT  4.510 1.965 4.630 2.140 ;
        RECT  4.025 1.965 4.510 2.085 ;
        RECT  4.360 1.055 4.480 1.845 ;
        RECT  3.930 1.055 4.360 1.175 ;
        RECT  4.190 0.670 4.310 0.935 ;
        RECT  4.080 1.295 4.200 1.845 ;
        RECT  3.800 1.725 4.080 1.845 ;
        RECT  3.930 0.370 4.060 0.540 ;
        RECT  3.905 1.965 4.025 2.140 ;
        RECT  3.810 0.370 3.930 1.590 ;
        RECT  1.610 2.020 3.905 2.140 ;
        RECT  3.775 1.330 3.810 1.590 ;
        RECT  3.680 1.725 3.800 1.900 ;
        RECT  2.000 1.780 3.680 1.900 ;
        RECT  3.510 0.830 3.630 1.615 ;
        RECT  3.340 0.830 3.510 0.950 ;
        RECT  3.480 1.495 3.510 1.615 ;
        RECT  3.360 1.495 3.480 1.660 ;
        RECT  2.240 1.540 3.360 1.660 ;
        RECT  3.170 0.445 3.340 0.950 ;
        RECT  2.875 0.780 3.170 0.950 ;
        RECT  2.640 1.300 2.880 1.420 ;
        RECT  2.840 0.830 2.875 0.950 ;
        RECT  2.695 0.400 2.865 0.590 ;
        RECT  2.640 0.420 2.695 0.590 ;
        RECT  2.520 0.420 2.640 1.420 ;
        RECT  1.650 0.420 2.520 0.540 ;
        RECT  2.000 0.660 2.400 0.780 ;
        RECT  2.120 1.330 2.240 1.660 ;
        RECT  1.880 0.660 2.000 1.900 ;
        RECT  1.640 0.750 1.760 1.830 ;
        RECT  1.530 0.420 1.650 0.630 ;
        RECT  1.500 0.750 1.640 0.870 ;
        RECT  1.545 1.400 1.640 1.830 ;
        RECT  1.490 1.950 1.610 2.140 ;
        RECT  0.955 0.510 1.530 0.630 ;
        RECT  0.635 1.950 1.490 2.070 ;
        RECT  0.955 1.025 1.475 1.195 ;
        RECT  0.835 0.420 0.955 1.825 ;
        RECT  0.785 0.420 0.835 0.850 ;
        RECT  0.785 1.395 0.835 1.825 ;
        RECT  0.515 0.465 0.635 2.070 ;
        RECT  0.445 0.465 0.515 0.895 ;
        RECT  0.445 1.640 0.515 2.070 ;
    END
END ACCSHCONX4AD
MACRO ACCSIHCONX2AD
    CLASS CORE ;
    FOREIGN ACCSIHCONX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 0.540 1.780 1.545 ;
        RECT  1.660 0.540 1.680 1.995 ;
        RECT  1.395 0.540 1.660 0.660 ;
        RECT  1.470 1.425 1.660 1.995 ;
        RECT  1.225 0.490 1.395 0.660 ;
        END
        AntennaDiffArea 0.396 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.520 1.605 0.690 2.050 ;
        RECT  0.210 1.605 0.520 1.725 ;
        RECT  0.240 0.410 0.410 0.840 ;
        RECT  0.210 0.720 0.240 0.840 ;
        RECT  0.070 0.720 0.210 1.725 ;
        END
        AntennaDiffArea 0.405 ;
    END CO0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.020 1.175 1.280 ;
        RECT  1.030 1.020 1.150 1.485 ;
        RECT  0.510 1.365 1.030 1.485 ;
        RECT  0.350 1.020 0.510 1.485 ;
        END
        AntennaGateArea 0.324 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.480 1.000 1.525 1.260 ;
        RECT  1.360 0.780 1.480 1.260 ;
        RECT  0.845 0.780 1.360 0.900 ;
        RECT  0.630 0.780 0.845 1.240 ;
        END
        AntennaGateArea 0.324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.760 -0.210 1.960 0.210 ;
        RECT  1.590 -0.210 1.760 0.415 ;
        RECT  1.010 -0.210 1.590 0.210 ;
        RECT  0.890 -0.210 1.010 0.580 ;
        RECT  0.000 -0.210 0.890 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 2.310 1.960 2.730 ;
        RECT  0.880 1.620 1.050 2.730 ;
        RECT  0.325 2.310 0.880 2.730 ;
        RECT  0.155 1.845 0.325 2.730 ;
        RECT  0.000 2.310 0.155 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
	 END
END ACCSIHCONX2AD
MACRO ACCSIHCONX4AD
    CLASS CORE ;
    FOREIGN ACCSIHCONX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.825 3.290 1.795 ;
        RECT  2.765 0.825 3.150 0.955 ;
        RECT  2.500 1.350 3.150 1.480 ;
        RECT  2.635 0.530 2.765 0.955 ;
        RECT  1.810 0.530 2.635 0.660 ;
        RECT  2.370 1.350 2.500 2.050 ;
        RECT  2.240 1.620 2.370 2.050 ;
        END
        AntennaDiffArea 0.63 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.255 1.570 1.425 2.030 ;
        RECT  0.690 1.570 1.255 1.700 ;
        RECT  1.030 0.615 1.055 0.745 ;
        RECT  0.910 0.485 1.030 0.745 ;
        RECT  0.210 0.615 0.910 0.745 ;
        RECT  0.520 1.570 0.690 2.030 ;
        RECT  0.210 1.570 0.520 1.700 ;
        RECT  0.070 0.615 0.210 1.700 ;
        END
        AntennaDiffArea 0.674 ;
    END CO0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 1.110 2.980 1.230 ;
        RECT  2.370 0.780 2.490 1.230 ;
        RECT  1.905 0.780 2.370 0.900 ;
        RECT  1.760 0.780 1.905 1.195 ;
        RECT  1.735 0.865 1.760 1.195 ;
        RECT  1.170 0.865 1.735 0.990 ;
        RECT  1.160 0.865 1.170 1.175 ;
        RECT  0.910 0.865 1.160 1.210 ;
        RECT  0.780 0.950 0.910 1.210 ;
        END
        AntennaGateArea 0.648 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.020 2.240 1.280 ;
        RECT  2.030 1.020 2.170 1.450 ;
        RECT  1.590 1.330 2.030 1.450 ;
        RECT  1.330 1.110 1.590 1.450 ;
        RECT  0.510 1.330 1.330 1.450 ;
        RECT  0.390 1.020 0.510 1.450 ;
        END
        AntennaGateArea 0.648 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.190 -0.210 3.360 0.210 ;
        RECT  2.930 -0.210 3.190 0.705 ;
        RECT  2.450 -0.210 2.930 0.210 ;
        RECT  2.190 -0.210 2.450 0.410 ;
        RECT  1.665 -0.210 2.190 0.210 ;
        RECT  1.495 -0.210 1.665 0.705 ;
        RECT  0.320 -0.210 1.495 0.210 ;
        RECT  0.150 -0.210 0.320 0.495 ;
        RECT  0.000 -0.210 0.150 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.030 2.310 3.360 2.730 ;
        RECT  2.850 1.600 3.030 2.730 ;
        RECT  1.785 2.310 2.850 2.730 ;
        RECT  1.615 1.600 1.785 2.730 ;
        RECT  1.060 2.310 1.615 2.730 ;
        RECT  0.890 1.845 1.060 2.730 ;
        RECT  0.325 2.310 0.890 2.730 ;
        RECT  0.155 1.845 0.325 2.730 ;
        RECT  0.000 2.310 0.155 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
	 END
END ACCSIHCONX4AD
MACRO ACHCINX2AD
    CLASS CORE ;
    FOREIGN ACHCINX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.150 0.870 5.270 1.850 ;
        RECT  4.745 0.870 5.150 0.990 ;
        RECT  4.950 1.690 5.150 1.850 ;
        RECT  4.520 1.690 4.950 1.810 ;
        RECT  4.485 0.350 4.745 0.990 ;
        RECT  4.400 1.690 4.520 2.140 ;
        RECT  4.125 2.020 4.400 2.140 ;
        END
        AntennaDiffArea 0.55 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.670 0.865 5.810 1.375 ;
        RECT  5.630 1.000 5.670 1.260 ;
        END
        AntennaGateArea 0.1613 ;
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 0.990 3.570 1.655 ;
        RECT  3.330 0.990 3.430 1.250 ;
        END
        AntennaGateArea 0.4086 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.000 0.350 1.260 ;
        RECT  0.070 1.000 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.510 -0.210 5.880 0.210 ;
        RECT  5.250 -0.210 5.510 0.500 ;
        RECT  3.765 -0.210 5.250 0.210 ;
        RECT  3.505 -0.210 3.765 0.320 ;
        RECT  0.730 -0.210 3.505 0.210 ;
        RECT  0.470 -0.210 0.730 0.260 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.460 2.310 5.880 2.730 ;
        RECT  5.200 2.210 5.460 2.730 ;
        RECT  3.640 2.310 5.200 2.730 ;
        RECT  3.380 2.020 3.640 2.730 ;
        RECT  0.615 2.310 3.380 2.730 ;
        RECT  0.445 1.800 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.880 2.520 ;
        LAYER M1 ;
        RECT  5.510 1.570 5.770 2.090 ;
        RECT  5.390 0.620 5.510 2.090 ;
        RECT  5.085 0.620 5.390 0.740 ;
        RECT  4.760 1.970 5.390 2.090 ;
        RECT  4.955 0.430 5.085 0.740 ;
        RECT  4.315 1.150 5.030 1.290 ;
        RECT  4.280 1.450 4.990 1.570 ;
        RECT  4.640 1.930 4.760 2.190 ;
        RECT  4.195 0.440 4.315 1.290 ;
        RECT  4.160 1.450 4.280 1.895 ;
        RECT  2.500 0.440 4.195 0.560 ;
        RECT  4.170 1.150 4.195 1.290 ;
        RECT  3.190 1.775 4.160 1.895 ;
        RECT  4.050 0.690 4.075 0.950 ;
        RECT  4.040 0.690 4.050 1.400 ;
        RECT  3.930 0.690 4.040 1.655 ;
        RECT  3.920 1.310 3.930 1.655 ;
        RECT  3.790 1.485 3.920 1.655 ;
        RECT  3.690 0.715 3.810 1.260 ;
        RECT  3.210 0.715 3.690 0.835 ;
        RECT  3.090 0.715 3.210 1.620 ;
        RECT  3.070 1.775 3.190 2.130 ;
        RECT  2.830 1.170 3.090 1.450 ;
        RECT  0.920 2.010 3.070 2.130 ;
        RECT  2.710 1.630 2.900 1.890 ;
        RECT  2.715 0.735 2.885 0.950 ;
        RECT  2.710 0.830 2.715 0.950 ;
        RECT  2.590 0.830 2.710 1.890 ;
        RECT  1.160 1.770 2.590 1.890 ;
        RECT  2.470 0.440 2.500 0.745 ;
        RECT  2.350 0.440 2.470 1.650 ;
        RECT  2.140 0.580 2.230 1.620 ;
        RECT  2.110 0.380 2.140 1.620 ;
        RECT  2.020 0.380 2.110 0.840 ;
        RECT  1.710 1.500 2.110 1.620 ;
        RECT  0.680 0.380 2.020 0.500 ;
        RECT  1.870 1.070 1.990 1.330 ;
        RECT  1.400 1.150 1.870 1.330 ;
        RECT  0.920 0.620 1.845 0.740 ;
        RECT  1.280 1.150 1.400 1.410 ;
        RECT  1.160 0.860 1.300 1.020 ;
        RECT  1.040 0.860 1.160 1.890 ;
        RECT  0.800 0.620 0.920 2.130 ;
        RECT  0.560 0.380 0.680 1.615 ;
        RECT  0.255 0.380 0.560 0.500 ;
        RECT  0.230 1.495 0.560 1.615 ;
        RECT  0.085 0.380 0.255 0.850 ;
        RECT  0.110 1.495 0.230 2.085 ;
    END
END ACHCINX2AD
MACRO ACHCINX4AD
    CLASS CORE ;
    FOREIGN ACHCINX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.955 0.645 6.105 1.720 ;
        RECT  5.950 0.645 5.955 1.350 ;
        RECT  5.275 0.645 5.950 0.770 ;
        RECT  5.505 1.220 5.950 1.350 ;
        RECT  5.375 1.220 5.505 2.125 ;
        RECT  4.915 2.005 5.375 2.125 ;
        RECT  5.105 0.340 5.275 0.770 ;
        END
        AntennaDiffArea 0.711 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.930 1.045 6.965 1.215 ;
        RECT  6.510 1.045 6.930 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.945 0.910 4.175 1.330 ;
        END
        AntennaGateArea 0.4718 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.000 0.350 1.260 ;
        RECT  0.070 1.000 0.210 1.375 ;
        END
        AntennaGateArea 0.1605 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.185 -0.210 7.280 0.210 ;
        RECT  7.015 -0.210 7.185 0.850 ;
        RECT  6.440 -0.210 7.015 0.210 ;
        RECT  6.180 -0.210 6.440 0.285 ;
        RECT  4.345 -0.210 6.180 0.210 ;
        RECT  4.085 -0.210 4.345 0.300 ;
        RECT  0.940 -0.210 4.085 0.210 ;
        RECT  0.420 -0.210 0.940 0.260 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.185 2.310 7.280 2.730 ;
        RECT  7.160 1.580 7.185 2.730 ;
        RECT  7.040 1.535 7.160 2.730 ;
        RECT  7.015 1.580 7.040 2.730 ;
        RECT  6.510 2.310 7.015 2.730 ;
        RECT  6.250 2.080 6.510 2.730 ;
        RECT  4.455 2.310 6.250 2.730 ;
        RECT  4.195 2.000 4.455 2.730 ;
        RECT  0.615 2.310 4.195 2.730 ;
        RECT  0.445 1.785 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.280 2.520 ;
        LAYER M1 ;
        RECT  6.655 0.420 6.825 0.850 ;
        RECT  6.680 1.535 6.800 2.055 ;
        RECT  6.375 1.535 6.680 1.655 ;
        RECT  6.375 0.730 6.655 0.850 ;
        RECT  6.255 0.405 6.375 1.960 ;
        RECT  5.455 0.405 6.255 0.525 ;
        RECT  5.745 1.840 6.255 1.960 ;
        RECT  5.485 0.890 5.745 1.050 ;
        RECT  5.625 1.540 5.745 2.060 ;
        RECT  4.955 0.890 5.485 1.010 ;
        RECT  5.135 1.130 5.255 1.880 ;
        RECT  4.075 1.760 5.135 1.880 ;
        RECT  4.835 0.420 4.955 1.400 ;
        RECT  3.260 0.420 4.835 0.540 ;
        RECT  4.715 1.520 4.815 1.640 ;
        RECT  4.595 0.680 4.715 1.640 ;
        RECT  4.555 1.520 4.595 1.640 ;
        RECT  4.355 0.660 4.475 1.270 ;
        RECT  3.805 0.660 4.355 0.780 ;
        RECT  3.805 1.520 4.095 1.640 ;
        RECT  3.955 1.760 4.075 2.140 ;
        RECT  0.855 2.020 3.955 2.140 ;
        RECT  3.685 0.660 3.805 1.640 ;
        RECT  3.565 1.780 3.755 1.900 ;
        RECT  3.445 0.660 3.685 0.780 ;
        RECT  3.445 0.930 3.565 1.900 ;
        RECT  3.020 0.930 3.445 1.050 ;
        RECT  1.160 1.780 3.445 1.900 ;
        RECT  3.205 1.170 3.325 1.660 ;
        RECT  3.140 0.385 3.260 0.810 ;
        RECT  2.540 1.170 3.205 1.290 ;
        RECT  2.540 0.385 3.140 0.505 ;
        RECT  2.300 1.415 3.035 1.535 ;
        RECT  2.900 0.670 3.020 1.050 ;
        RECT  2.710 0.670 2.900 0.790 ;
        RECT  2.420 0.385 2.540 1.290 ;
        RECT  2.180 0.880 2.300 1.660 ;
        RECT  2.160 0.880 2.180 1.000 ;
        RECT  1.680 1.540 2.180 1.660 ;
        RECT  2.040 0.380 2.160 1.000 ;
        RECT  0.680 0.380 2.040 0.500 ;
        RECT  1.885 1.150 2.005 1.410 ;
        RECT  1.400 1.290 1.885 1.410 ;
        RECT  1.650 0.620 1.820 0.790 ;
        RECT  0.920 0.620 1.650 0.740 ;
        RECT  1.160 0.870 1.505 0.990 ;
        RECT  1.280 1.290 1.400 1.605 ;
        RECT  1.040 0.870 1.160 1.900 ;
        RECT  0.975 1.640 1.040 1.900 ;
        RECT  0.855 0.620 0.920 1.500 ;
        RECT  0.800 0.620 0.855 2.140 ;
        RECT  0.735 1.380 0.800 2.140 ;
        RECT  0.590 0.380 0.680 1.260 ;
        RECT  0.560 0.380 0.590 1.615 ;
        RECT  0.255 0.380 0.560 0.500 ;
        RECT  0.470 1.000 0.560 1.615 ;
        RECT  0.255 1.495 0.470 1.615 ;
        RECT  0.085 0.380 0.255 0.810 ;
        RECT  0.100 1.495 0.255 2.085 ;
    END
END ACHCINX4AD
MACRO ACHCONX2AD
    CLASS CORE ;
    FOREIGN ACHCONX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.150 0.870 5.270 1.850 ;
        RECT  4.745 0.870 5.150 0.990 ;
        RECT  4.950 1.690 5.150 1.850 ;
        RECT  4.520 1.690 4.950 1.810 ;
        RECT  4.485 0.350 4.745 0.990 ;
        RECT  4.400 1.690 4.520 2.140 ;
        RECT  4.125 2.020 4.400 2.140 ;
        END
        AntennaDiffArea 0.55 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.670 0.865 5.810 1.375 ;
        RECT  5.630 1.000 5.670 1.260 ;
        END
        AntennaGateArea 0.1613 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.570 1.000 3.730 1.260 ;
        RECT  3.430 1.000 3.570 1.655 ;
        RECT  3.330 1.000 3.430 1.260 ;
        END
        AntennaGateArea 0.5621 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.000 0.350 1.260 ;
        RECT  0.070 1.000 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.510 -0.210 5.880 0.210 ;
        RECT  5.250 -0.210 5.510 0.500 ;
        RECT  3.765 -0.210 5.250 0.210 ;
        RECT  3.505 -0.210 3.765 0.320 ;
        RECT  0.730 -0.210 3.505 0.210 ;
        RECT  0.470 -0.210 0.730 0.260 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.460 2.310 5.880 2.730 ;
        RECT  5.200 2.210 5.460 2.730 ;
        RECT  3.640 2.310 5.200 2.730 ;
        RECT  3.380 2.020 3.640 2.730 ;
        RECT  0.615 2.310 3.380 2.730 ;
        RECT  0.445 1.800 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.880 2.520 ;
        LAYER M1 ;
        RECT  5.510 1.570 5.770 2.090 ;
        RECT  5.390 0.620 5.510 2.090 ;
        RECT  5.085 0.620 5.390 0.740 ;
        RECT  4.760 1.970 5.390 2.090 ;
        RECT  4.955 0.430 5.085 0.740 ;
        RECT  4.315 1.150 5.030 1.290 ;
        RECT  4.280 1.450 4.990 1.570 ;
        RECT  4.640 1.930 4.760 2.190 ;
        RECT  4.195 0.440 4.315 1.290 ;
        RECT  4.160 1.450 4.280 1.895 ;
        RECT  2.500 0.440 4.195 0.560 ;
        RECT  4.170 1.150 4.195 1.290 ;
        RECT  3.190 1.775 4.160 1.895 ;
        RECT  4.040 0.690 4.075 0.950 ;
        RECT  3.920 0.690 4.040 1.655 ;
        RECT  3.790 1.485 3.920 1.655 ;
        RECT  3.210 0.715 3.375 0.835 ;
        RECT  3.090 0.715 3.210 1.620 ;
        RECT  3.070 1.775 3.190 2.130 ;
        RECT  2.830 1.170 3.090 1.450 ;
        RECT  0.920 2.010 3.070 2.130 ;
        RECT  2.710 1.630 2.900 1.890 ;
        RECT  2.715 0.735 2.885 0.950 ;
        RECT  2.710 0.830 2.715 0.950 ;
        RECT  2.590 0.830 2.710 1.890 ;
        RECT  1.160 1.770 2.590 1.890 ;
        RECT  2.470 0.440 2.500 0.745 ;
        RECT  2.350 0.440 2.470 1.650 ;
        RECT  2.140 0.580 2.230 1.620 ;
        RECT  2.110 0.380 2.140 1.620 ;
        RECT  2.020 0.380 2.110 0.840 ;
        RECT  1.710 1.500 2.110 1.620 ;
        RECT  0.680 0.380 2.020 0.500 ;
        RECT  1.870 1.070 1.990 1.330 ;
        RECT  1.400 1.150 1.870 1.330 ;
        RECT  0.920 0.620 1.845 0.740 ;
        RECT  1.280 1.150 1.400 1.410 ;
        RECT  1.160 0.860 1.300 1.020 ;
        RECT  1.040 0.860 1.160 1.890 ;
        RECT  0.800 0.620 0.920 2.130 ;
        RECT  0.560 0.380 0.680 1.615 ;
        RECT  0.255 0.380 0.560 0.500 ;
        RECT  0.230 1.495 0.560 1.615 ;
        RECT  0.085 0.380 0.255 0.850 ;
        RECT  0.110 1.495 0.230 2.085 ;
    END
END ACHCONX2AD
MACRO ACHCONX4AD
    CLASS CORE ;
    FOREIGN ACHCONX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.955 0.645 6.105 1.720 ;
        RECT  5.950 0.645 5.955 1.350 ;
        RECT  5.275 0.645 5.950 0.770 ;
        RECT  5.505 1.220 5.950 1.350 ;
        RECT  5.375 1.220 5.505 2.125 ;
        RECT  4.915 2.005 5.375 2.125 ;
        RECT  5.105 0.340 5.275 0.770 ;
        END
        AntennaDiffArea 0.711 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.930 1.045 6.965 1.215 ;
        RECT  6.510 1.045 6.930 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.945 0.910 4.420 1.225 ;
        END
        AntennaGateArea 0.5953 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.000 0.350 1.260 ;
        RECT  0.070 1.000 0.210 1.375 ;
        END
        AntennaGateArea 0.1605 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.185 -0.210 7.280 0.210 ;
        RECT  7.015 -0.210 7.185 0.850 ;
        RECT  6.440 -0.210 7.015 0.210 ;
        RECT  6.180 -0.210 6.440 0.285 ;
        RECT  4.345 -0.210 6.180 0.210 ;
        RECT  4.085 -0.210 4.345 0.300 ;
        RECT  0.940 -0.210 4.085 0.210 ;
        RECT  0.420 -0.210 0.940 0.260 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.185 2.310 7.280 2.730 ;
        RECT  7.160 1.580 7.185 2.730 ;
        RECT  7.040 1.535 7.160 2.730 ;
        RECT  7.015 1.580 7.040 2.730 ;
        RECT  6.510 2.310 7.015 2.730 ;
        RECT  6.250 2.080 6.510 2.730 ;
        RECT  4.455 2.310 6.250 2.730 ;
        RECT  4.195 2.000 4.455 2.730 ;
        RECT  0.615 2.310 4.195 2.730 ;
        RECT  0.445 1.785 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.280 2.520 ;
        LAYER M1 ;
        RECT  6.655 0.420 6.825 0.850 ;
        RECT  6.680 1.535 6.800 2.055 ;
        RECT  6.375 1.535 6.680 1.655 ;
        RECT  6.375 0.730 6.655 0.850 ;
        RECT  6.255 0.405 6.375 1.960 ;
        RECT  5.455 0.405 6.255 0.525 ;
        RECT  5.745 1.840 6.255 1.960 ;
        RECT  5.485 0.890 5.745 1.050 ;
        RECT  5.625 1.540 5.745 2.060 ;
        RECT  4.955 0.890 5.485 1.010 ;
        RECT  5.135 1.130 5.255 1.880 ;
        RECT  4.075 1.760 5.135 1.880 ;
        RECT  4.835 0.420 4.955 1.400 ;
        RECT  3.260 0.420 4.835 0.540 ;
        RECT  4.715 1.520 4.815 1.640 ;
        RECT  4.595 0.680 4.715 1.640 ;
        RECT  4.555 1.520 4.595 1.640 ;
        RECT  3.805 1.520 4.095 1.640 ;
        RECT  3.955 1.760 4.075 2.140 ;
        RECT  3.805 0.660 3.965 0.780 ;
        RECT  0.855 2.020 3.955 2.140 ;
        RECT  3.685 0.660 3.805 1.640 ;
        RECT  3.565 1.780 3.755 1.900 ;
        RECT  3.445 0.660 3.685 0.780 ;
        RECT  3.445 0.930 3.565 1.900 ;
        RECT  3.020 0.930 3.445 1.050 ;
        RECT  1.160 1.780 3.445 1.900 ;
        RECT  3.205 1.170 3.325 1.660 ;
        RECT  3.140 0.385 3.260 0.810 ;
        RECT  2.540 1.170 3.205 1.290 ;
        RECT  2.540 0.385 3.140 0.505 ;
        RECT  2.300 1.415 3.035 1.535 ;
        RECT  2.900 0.670 3.020 1.050 ;
        RECT  2.710 0.670 2.900 0.790 ;
        RECT  2.420 0.385 2.540 1.290 ;
        RECT  2.180 0.880 2.300 1.660 ;
        RECT  2.160 0.880 2.180 1.000 ;
        RECT  1.680 1.540 2.180 1.660 ;
        RECT  2.040 0.380 2.160 1.000 ;
        RECT  0.680 0.380 2.040 0.500 ;
        RECT  1.885 1.150 2.005 1.410 ;
        RECT  1.400 1.290 1.885 1.410 ;
        RECT  1.650 0.620 1.820 0.790 ;
        RECT  0.920 0.620 1.650 0.740 ;
        RECT  1.160 0.870 1.505 0.990 ;
        RECT  1.280 1.290 1.400 1.605 ;
        RECT  1.040 0.870 1.160 1.900 ;
        RECT  0.975 1.640 1.040 1.900 ;
        RECT  0.855 0.620 0.920 1.500 ;
        RECT  0.800 0.620 0.855 2.140 ;
        RECT  0.735 1.380 0.800 2.140 ;
        RECT  0.590 0.380 0.680 1.260 ;
        RECT  0.560 0.380 0.590 1.615 ;
        RECT  0.255 0.380 0.560 0.500 ;
        RECT  0.470 1.000 0.560 1.615 ;
        RECT  0.255 1.495 0.470 1.615 ;
        RECT  0.085 0.380 0.255 0.810 ;
        RECT  0.100 1.495 0.255 2.085 ;
    END
END ACHCONX4AD
MACRO ADDFHX1AD
    CLASS CORE ;
    FOREIGN ADDFHX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.035 0.690 8.050 1.555 ;
        RECT  7.910 0.690 8.035 1.840 ;
        RECT  7.865 0.690 7.910 0.860 ;
        RECT  7.865 1.410 7.910 1.840 ;
        END
        AntennaDiffArea 0.203 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.350 0.700 7.490 1.620 ;
        RECT  7.120 0.700 7.350 0.870 ;
        RECT  7.120 1.450 7.350 1.620 ;
        END
        AntennaDiffArea 0.204 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.720 0.865 6.930 1.375 ;
        END
        AntennaGateArea 0.0994 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.520 0.860 3.640 1.380 ;
        RECT  3.385 1.190 3.520 1.380 ;
        END
        AntennaGateArea 0.379 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 1.010 0.360 1.270 ;
        RECT  0.070 0.865 0.240 1.375 ;
        END
        AntennaGateArea 0.1618 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.655 -0.210 8.120 0.210 ;
        RECT  7.485 -0.210 7.655 0.385 ;
        RECT  6.680 -0.210 7.485 0.210 ;
        RECT  6.420 -0.210 6.680 0.320 ;
        RECT  4.450 -0.210 6.420 0.210 ;
        RECT  4.190 -0.210 4.450 0.300 ;
        RECT  1.025 -0.210 4.190 0.210 ;
        RECT  0.505 -0.210 1.025 0.320 ;
        RECT  0.000 -0.210 0.505 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.725 2.310 8.120 2.730 ;
        RECT  7.465 2.220 7.725 2.730 ;
        RECT  6.615 2.310 7.465 2.730 ;
        RECT  6.355 2.220 6.615 2.730 ;
        RECT  4.080 2.310 6.355 2.730 ;
        RECT  3.960 1.950 4.080 2.730 ;
        RECT  0.970 2.310 3.960 2.730 ;
        RECT  0.970 1.940 1.055 2.110 ;
        RECT  0.710 1.940 0.970 2.730 ;
        RECT  0.625 1.940 0.710 2.110 ;
        RECT  0.000 2.310 0.710 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.120 2.520 ;
        LAYER M1 ;
        RECT  7.730 1.010 7.770 1.270 ;
        RECT  7.610 1.010 7.730 1.860 ;
        RECT  5.860 1.740 7.610 1.860 ;
        RECT  7.085 1.980 7.345 2.190 ;
        RECT  5.110 1.980 7.085 2.100 ;
        RECT  6.800 0.380 7.060 0.560 ;
        RECT  6.490 1.500 6.995 1.620 ;
        RECT  6.490 0.440 6.800 0.560 ;
        RECT  6.350 0.440 6.490 1.620 ;
        RECT  5.570 0.440 6.350 0.560 ;
        RECT  6.100 0.680 6.230 1.585 ;
        RECT  6.060 1.415 6.100 1.585 ;
        RECT  5.740 0.680 5.860 1.860 ;
        RECT  5.625 1.740 5.740 1.860 ;
        RECT  5.450 0.440 5.570 0.895 ;
        RECT  5.430 1.685 5.480 1.855 ;
        RECT  5.430 0.725 5.450 0.895 ;
        RECT  5.310 0.725 5.430 1.855 ;
        RECT  5.070 0.360 5.330 0.540 ;
        RECT  5.110 0.725 5.165 0.895 ;
        RECT  4.990 0.725 5.110 2.190 ;
        RECT  4.200 0.420 5.070 0.540 ;
        RECT  4.640 2.070 4.990 2.190 ;
        RECT  4.750 0.660 4.870 1.950 ;
        RECT  4.570 0.660 4.750 0.780 ;
        RECT  4.465 1.830 4.750 1.950 ;
        RECT  4.460 0.900 4.630 1.710 ;
        RECT  4.320 1.830 4.465 2.065 ;
        RECT  4.200 0.900 4.460 1.100 ;
        RECT  4.200 1.710 4.320 2.065 ;
        RECT  3.880 1.260 4.315 1.440 ;
        RECT  4.090 0.420 4.200 1.100 ;
        RECT  3.460 1.710 4.200 1.830 ;
        RECT  4.000 0.380 4.090 1.100 ;
        RECT  2.740 0.380 4.000 0.500 ;
        RECT  3.760 0.620 3.880 1.440 ;
        RECT  2.980 0.620 3.760 0.740 ;
        RECT  3.340 1.500 3.460 2.020 ;
        RECT  3.220 0.860 3.400 0.980 ;
        RECT  3.100 0.860 3.220 2.140 ;
        RECT  1.540 2.020 3.100 2.140 ;
        RECT  2.860 0.620 2.980 1.900 ;
        RECT  1.900 1.780 2.860 1.900 ;
        RECT  2.620 0.380 2.740 1.660 ;
        RECT  2.430 1.540 2.620 1.660 ;
        RECT  2.330 0.505 2.500 0.765 ;
        RECT  2.290 0.380 2.330 0.765 ;
        RECT  2.170 0.380 2.290 1.660 ;
        RECT  1.250 0.380 2.170 0.500 ;
        RECT  2.115 1.490 2.170 1.660 ;
        RECT  1.900 0.630 2.050 0.800 ;
        RECT  1.780 0.630 1.900 1.900 ;
        RECT  1.540 0.630 1.565 0.800 ;
        RECT  1.395 0.630 1.540 2.140 ;
        RECT  1.130 0.380 1.250 0.560 ;
        RECT  0.925 1.085 1.205 1.345 ;
        RECT  0.610 0.440 1.130 0.560 ;
        RECT  0.755 0.735 0.925 1.585 ;
        RECT  0.490 0.440 0.610 1.615 ;
        RECT  0.085 0.575 0.490 0.745 ;
        RECT  0.255 1.495 0.490 1.615 ;
        RECT  0.085 1.495 0.255 1.925 ;
    END
END ADDFHX1AD
MACRO ADDFHX2AD
    CLASS CORE ;
    FOREIGN ADDFHX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.835 0.800 10.850 1.500 ;
        RECT  10.820 0.410 10.835 1.500 ;
        RECT  10.710 0.410 10.820 2.025 ;
        RECT  10.695 0.410 10.710 0.940 ;
        RECT  10.680 1.360 10.710 2.025 ;
        RECT  10.665 0.410 10.695 0.840 ;
        END
        AntennaDiffArea 0.373 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.115 0.865 10.290 1.375 ;
        RECT  9.995 0.735 10.115 1.620 ;
        RECT  9.945 0.735 9.995 0.905 ;
        RECT  9.945 1.450 9.995 1.620 ;
        END
        AntennaDiffArea 0.315 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.565 0.865 9.775 1.375 ;
        END
        AntennaGateArea 0.1605 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.185 1.190 6.635 1.450 ;
        END
        AntennaGateArea 0.6782 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.060 0.695 1.230 ;
        RECT  0.070 0.865 0.210 1.655 ;
        END
        AntennaGateArea 0.2872 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.475 -0.210 10.920 0.210 ;
        RECT  10.305 -0.210 10.475 0.745 ;
        RECT  9.500 -0.210 10.305 0.210 ;
        RECT  9.240 -0.210 9.500 0.290 ;
        RECT  6.595 -0.210 9.240 0.210 ;
        RECT  6.425 -0.210 6.595 0.255 ;
        RECT  1.890 -0.210 6.425 0.210 ;
        RECT  1.720 -0.210 1.890 0.255 ;
        RECT  0.855 -0.210 1.720 0.210 ;
        RECT  0.165 -0.210 0.855 0.255 ;
        RECT  0.000 -0.210 0.165 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.475 2.310 10.920 2.730 ;
        RECT  10.305 1.980 10.475 2.730 ;
        RECT  9.345 2.310 10.305 2.730 ;
        RECT  9.085 2.220 9.345 2.730 ;
        RECT  6.500 2.310 9.085 2.730 ;
        RECT  6.330 1.870 6.500 2.730 ;
        RECT  1.755 2.310 6.330 2.730 ;
        RECT  1.585 2.025 1.755 2.730 ;
        RECT  0.880 2.310 1.585 2.730 ;
        RECT  0.100 2.230 0.880 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.920 2.520 ;
        LAYER M1 ;
        RECT  10.545 1.020 10.590 1.280 ;
        RECT  10.425 1.020 10.545 1.860 ;
        RECT  8.535 1.740 10.425 1.860 ;
        RECT  9.710 1.980 9.970 2.185 ;
        RECT  9.665 0.360 9.835 0.530 ;
        RECT  9.260 1.500 9.805 1.620 ;
        RECT  8.580 1.980 9.710 2.100 ;
        RECT  9.445 0.410 9.665 0.530 ;
        RECT  9.325 0.410 9.445 1.040 ;
        RECT  8.400 0.410 9.325 0.530 ;
        RECT  9.260 0.920 9.325 1.040 ;
        RECT  9.140 0.920 9.260 1.620 ;
        RECT  9.050 1.025 9.140 1.285 ;
        RECT  8.930 0.680 9.120 0.800 ;
        RECT  8.930 1.500 8.965 1.620 ;
        RECT  8.810 0.680 8.930 1.620 ;
        RECT  8.705 1.500 8.810 1.620 ;
        RECT  8.570 0.650 8.690 1.000 ;
        RECT  8.490 1.980 8.580 2.125 ;
        RECT  8.535 0.880 8.570 1.000 ;
        RECT  8.415 0.880 8.535 1.860 ;
        RECT  7.935 2.005 8.490 2.125 ;
        RECT  8.295 0.410 8.400 0.755 ;
        RECT  8.280 0.410 8.295 1.880 ;
        RECT  8.175 0.585 8.280 1.880 ;
        RECT  8.055 1.620 8.175 1.880 ;
        RECT  7.935 0.585 7.970 0.845 ;
        RECT  7.815 0.585 7.935 2.125 ;
        RECT  7.070 1.850 7.815 1.980 ;
        RECT  7.575 0.585 7.695 1.730 ;
        RECT  7.490 0.585 7.575 0.845 ;
        RECT  6.860 1.610 7.575 1.730 ;
        RECT  7.250 0.335 7.370 1.410 ;
        RECT  7.110 0.335 7.250 0.540 ;
        RECT  6.885 1.290 7.250 1.410 ;
        RECT  7.010 0.665 7.130 1.150 ;
        RECT  6.280 0.420 7.110 0.540 ;
        RECT  6.070 0.665 7.010 0.785 ;
        RECT  6.715 0.905 6.885 1.075 ;
        RECT  6.690 1.610 6.860 2.060 ;
        RECT  6.025 0.905 6.715 1.025 ;
        RECT  6.140 1.610 6.690 1.730 ;
        RECT  6.160 0.380 6.280 0.540 ;
        RECT  5.015 0.380 6.160 0.500 ;
        RECT  6.025 1.610 6.140 2.060 ;
        RECT  5.950 0.620 6.070 0.785 ;
        RECT  5.905 0.905 6.025 2.060 ;
        RECT  5.255 0.620 5.950 0.740 ;
        RECT  5.665 1.000 5.785 2.140 ;
        RECT  5.545 1.000 5.665 1.120 ;
        RECT  2.090 2.020 5.665 2.140 ;
        RECT  5.375 0.860 5.545 1.120 ;
        RECT  5.425 1.240 5.545 1.900 ;
        RECT  5.255 1.240 5.425 1.360 ;
        RECT  2.635 1.780 5.425 1.900 ;
        RECT  5.015 1.540 5.305 1.660 ;
        RECT  5.135 0.620 5.255 1.360 ;
        RECT  4.930 0.380 5.015 1.660 ;
        RECT  4.895 0.365 4.930 1.660 ;
        RECT  4.855 0.365 4.895 0.500 ;
        RECT  4.015 1.540 4.895 1.660 ;
        RECT  4.480 0.365 4.855 0.485 ;
        RECT  4.710 0.605 4.760 0.775 ;
        RECT  4.590 0.605 4.710 1.420 ;
        RECT  3.895 1.300 4.590 1.420 ;
        RECT  4.410 0.365 4.480 0.500 ;
        RECT  4.400 0.380 4.410 0.500 ;
        RECT  4.230 0.380 4.400 0.660 ;
        RECT  3.895 0.385 4.040 0.725 ;
        RECT  3.775 0.385 3.895 1.610 ;
        RECT  2.130 0.385 3.775 0.505 ;
        RECT  3.160 1.490 3.775 1.610 ;
        RECT  3.535 0.625 3.655 1.225 ;
        RECT  2.695 1.105 3.535 1.225 ;
        RECT  2.900 1.490 3.160 1.660 ;
        RECT  2.885 0.625 3.005 0.950 ;
        RECT  2.325 0.625 2.885 0.745 ;
        RECT  2.635 0.865 2.695 1.225 ;
        RECT  2.515 0.865 2.635 1.900 ;
        RECT  2.435 0.865 2.515 0.985 ;
        RECT  2.305 1.655 2.515 1.900 ;
        RECT  2.220 0.625 2.325 0.800 ;
        RECT  2.090 0.680 2.220 0.800 ;
        RECT  2.035 0.385 2.130 0.540 ;
        RECT  1.970 0.680 2.090 2.140 ;
        RECT  0.935 0.420 2.035 0.540 ;
        RECT  1.360 0.680 1.970 0.800 ;
        RECT  1.440 1.705 1.970 1.825 ;
        RECT  1.235 1.105 1.850 1.275 ;
        RECT  1.320 1.705 1.440 2.140 ;
        RECT  1.180 2.020 1.320 2.140 ;
        RECT  1.065 0.690 1.235 1.585 ;
        RECT  0.815 0.420 0.935 1.605 ;
        RECT  0.385 0.675 0.815 0.845 ;
        RECT  0.555 1.435 0.815 1.605 ;
        RECT  0.385 1.435 0.555 1.865 ;
    END
END ADDFHX2AD
MACRO ADDFHX4AD
    CLASS CORE ;
    FOREIGN ADDFHX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  17.195 0.690 17.290 1.515 ;
        RECT  17.150 0.690 17.195 1.915 ;
        RECT  17.100 0.690 17.150 0.830 ;
        RECT  17.025 1.375 17.150 1.915 ;
        RECT  16.930 0.400 17.100 0.830 ;
        END
        AntennaDiffArea 0.422 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.450 1.395 16.475 1.565 ;
        RECT  16.210 0.440 16.450 1.565 ;
        END
        AntennaDiffArea 0.422 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  15.145 0.910 15.375 1.260 ;
        RECT  14.945 1.000 15.145 1.260 ;
        END
        AntennaGateArea 0.3226 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.610 1.145 8.750 1.305 ;
        RECT  8.190 1.145 8.610 1.375 ;
        END
        AntennaGateArea 1.2832 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.585 1.085 1.095 1.330 ;
        RECT  0.315 1.085 0.585 1.240 ;
        END
        AntennaGateArea 0.5745 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  17.530 -0.210 17.640 0.210 ;
        RECT  17.410 -0.210 17.530 0.880 ;
        RECT  16.740 -0.210 17.410 0.210 ;
        RECT  16.570 -0.210 16.740 0.830 ;
        RECT  16.020 -0.210 16.570 0.210 ;
        RECT  15.850 -0.210 16.020 0.830 ;
        RECT  15.320 -0.210 15.850 0.210 ;
        RECT  15.150 -0.210 15.320 0.435 ;
        RECT  14.275 -0.210 15.150 0.210 ;
        RECT  14.015 -0.210 14.275 0.260 ;
        RECT  9.415 -0.210 14.015 0.210 ;
        RECT  9.155 -0.210 9.415 0.260 ;
        RECT  8.585 -0.210 9.155 0.210 ;
        RECT  8.325 -0.210 8.585 0.260 ;
        RECT  2.820 -0.210 8.325 0.210 ;
        RECT  2.560 -0.210 2.820 0.300 ;
        RECT  2.060 -0.210 2.560 0.210 ;
        RECT  1.800 -0.210 2.060 0.300 ;
        RECT  1.400 -0.210 1.800 0.210 ;
        RECT  1.140 -0.210 1.400 0.300 ;
        RECT  0.615 -0.210 1.140 0.210 ;
        RECT  0.445 -0.210 0.615 0.680 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  17.555 2.310 17.640 2.730 ;
        RECT  17.385 1.680 17.555 2.730 ;
        RECT  16.835 2.310 17.385 2.730 ;
        RECT  16.665 2.040 16.835 2.730 ;
        RECT  16.090 2.310 16.665 2.730 ;
        RECT  15.970 1.985 16.090 2.730 ;
        RECT  15.220 2.310 15.970 2.730 ;
        RECT  14.960 2.220 15.220 2.730 ;
        RECT  14.100 2.310 14.960 2.730 ;
        RECT  13.840 2.220 14.100 2.730 ;
        RECT  9.285 2.310 13.840 2.730 ;
        RECT  9.115 1.940 9.285 2.730 ;
        RECT  8.565 2.310 9.115 2.730 ;
        RECT  8.395 1.880 8.565 2.730 ;
        RECT  2.755 2.310 8.395 2.730 ;
        RECT  2.585 1.770 2.755 2.730 ;
        RECT  2.035 2.310 2.585 2.730 ;
        RECT  1.865 1.490 2.035 2.730 ;
        RECT  1.335 2.310 1.865 2.730 ;
        RECT  1.165 1.715 1.335 2.730 ;
        RECT  0.615 2.310 1.165 2.730 ;
        RECT  0.445 1.715 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 17.640 2.520 ;
        LAYER M1 ;
        RECT  16.840 1.045 16.980 1.215 ;
        RECT  16.720 1.045 16.840 1.805 ;
        RECT  14.980 1.685 16.720 1.805 ;
        RECT  15.710 1.930 15.830 2.190 ;
        RECT  13.490 1.980 15.710 2.100 ;
        RECT  15.535 0.430 15.655 0.950 ;
        RECT  14.825 1.445 15.600 1.565 ;
        RECT  14.960 0.650 15.535 0.770 ;
        RECT  14.860 1.685 14.980 1.860 ;
        RECT  14.825 0.380 14.960 0.810 ;
        RECT  13.280 1.740 14.860 1.860 ;
        RECT  14.705 0.380 14.825 1.565 ;
        RECT  12.075 0.380 14.705 0.500 ;
        RECT  14.625 1.120 14.705 1.565 ;
        RECT  13.940 1.120 14.625 1.290 ;
        RECT  14.465 0.680 14.585 0.940 ;
        RECT  13.755 1.500 14.480 1.620 ;
        RECT  13.755 0.680 14.465 0.800 ;
        RECT  13.635 0.680 13.755 1.620 ;
        RECT  13.155 0.965 13.635 1.085 ;
        RECT  12.920 1.500 13.635 1.620 ;
        RECT  13.320 0.620 13.490 0.830 ;
        RECT  13.370 1.980 13.490 2.140 ;
        RECT  11.225 2.020 13.370 2.140 ;
        RECT  12.540 0.620 13.320 0.740 ;
        RECT  13.160 1.740 13.280 1.900 ;
        RECT  12.540 1.780 13.160 1.900 ;
        RECT  12.895 0.860 13.155 1.085 ;
        RECT  12.660 1.500 12.920 1.660 ;
        RECT  12.420 0.620 12.540 1.900 ;
        RECT  12.290 0.660 12.420 0.830 ;
        RECT  11.730 1.780 12.420 1.900 ;
        RECT  12.180 1.400 12.300 1.660 ;
        RECT  12.075 1.400 12.180 1.625 ;
        RECT  11.955 0.380 12.075 1.625 ;
        RECT  11.450 0.380 11.955 0.500 ;
        RECT  11.585 1.505 11.955 1.625 ;
        RECT  11.690 0.620 11.740 0.790 ;
        RECT  11.570 0.620 11.690 1.020 ;
        RECT  11.415 1.505 11.585 1.865 ;
        RECT  10.655 0.895 11.570 1.020 ;
        RECT  11.330 0.380 11.450 0.745 ;
        RECT  10.840 1.505 11.415 1.625 ;
        RECT  11.165 0.625 11.330 0.745 ;
        RECT  11.055 1.745 11.225 2.140 ;
        RECT  11.020 0.330 11.190 0.500 ;
        RECT  10.590 2.020 11.055 2.140 ;
        RECT  10.275 0.620 11.045 0.740 ;
        RECT  9.690 0.380 11.020 0.500 ;
        RECT  10.720 1.505 10.840 1.875 ;
        RECT  10.590 0.860 10.655 1.020 ;
        RECT  10.470 0.860 10.590 2.140 ;
        RECT  10.395 0.860 10.470 0.980 ;
        RECT  10.050 2.020 10.470 2.140 ;
        RECT  10.275 1.095 10.340 1.900 ;
        RECT  10.220 0.620 10.275 1.900 ;
        RECT  10.155 0.620 10.220 1.215 ;
        RECT  9.645 1.700 10.220 1.820 ;
        RECT  9.810 0.620 10.155 0.740 ;
        RECT  10.035 1.320 10.095 1.580 ;
        RECT  9.790 1.965 10.050 2.140 ;
        RECT  9.975 0.860 10.035 1.580 ;
        RECT  9.915 0.860 9.975 1.555 ;
        RECT  9.690 0.860 9.915 0.980 ;
        RECT  9.765 1.105 9.795 1.275 ;
        RECT  9.365 1.105 9.765 1.290 ;
        RECT  9.570 0.380 9.690 0.980 ;
        RECT  9.475 1.700 9.645 2.130 ;
        RECT  6.400 0.380 9.570 0.500 ;
        RECT  9.125 1.700 9.475 1.820 ;
        RECT  9.245 0.620 9.365 1.290 ;
        RECT  6.640 0.620 9.245 0.740 ;
        RECT  9.005 0.860 9.125 1.820 ;
        RECT  7.945 0.860 9.005 0.980 ;
        RECT  8.925 1.640 9.005 1.820 ;
        RECT  8.755 1.640 8.925 2.070 ;
        RECT  8.205 1.640 8.755 1.760 ;
        RECT  8.035 1.640 8.205 2.115 ;
        RECT  7.950 1.640 8.035 1.760 ;
        RECT  7.830 1.135 7.950 1.760 ;
        RECT  7.710 0.860 7.825 0.980 ;
        RECT  7.590 0.860 7.710 2.140 ;
        RECT  6.765 0.860 7.590 0.980 ;
        RECT  3.835 2.020 7.590 2.140 ;
        RECT  7.350 1.205 7.470 1.900 ;
        RECT  6.640 1.205 7.350 1.325 ;
        RECT  4.915 1.780 7.350 1.900 ;
        RECT  6.400 1.540 7.230 1.660 ;
        RECT  6.520 0.620 6.640 1.325 ;
        RECT  6.280 0.380 6.400 1.660 ;
        RECT  5.755 0.380 6.280 0.500 ;
        RECT  5.420 1.540 6.280 1.660 ;
        RECT  6.020 0.650 6.160 0.770 ;
        RECT  6.020 1.300 6.060 1.420 ;
        RECT  5.900 0.650 6.020 1.420 ;
        RECT  5.800 1.210 5.900 1.420 ;
        RECT  5.370 1.210 5.800 1.330 ;
        RECT  5.585 0.380 5.755 0.670 ;
        RECT  5.275 0.390 5.370 1.330 ;
        RECT  5.250 0.390 5.275 1.640 ;
        RECT  4.675 0.390 5.250 0.510 ;
        RECT  5.105 1.210 5.250 1.640 ;
        RECT  4.555 1.210 5.105 1.330 ;
        RECT  4.865 0.630 5.035 1.085 ;
        RECT  4.745 1.650 4.915 1.900 ;
        RECT  4.305 0.965 4.865 1.085 ;
        RECT  4.170 1.780 4.745 1.900 ;
        RECT  4.505 0.390 4.675 0.810 ;
        RECT  4.385 1.210 4.555 1.660 ;
        RECT  3.200 0.390 4.505 0.510 ;
        RECT  4.135 0.630 4.305 1.085 ;
        RECT  4.050 1.365 4.170 1.900 ;
        RECT  3.590 0.965 4.135 1.085 ;
        RECT  3.475 1.365 4.050 1.495 ;
        RECT  3.765 0.660 3.935 0.830 ;
        RECT  3.665 1.630 3.835 2.140 ;
        RECT  3.115 0.660 3.765 0.780 ;
        RECT  3.115 2.020 3.665 2.140 ;
        RECT  3.475 0.900 3.590 1.085 ;
        RECT  3.330 0.900 3.475 1.885 ;
        RECT  3.305 1.715 3.330 1.885 ;
        RECT  3.080 0.390 3.200 0.540 ;
        RECT  2.960 0.660 3.115 2.140 ;
        RECT  1.355 0.420 3.080 0.540 ;
        RECT  2.225 0.660 2.960 0.830 ;
        RECT  2.945 1.480 2.960 2.140 ;
        RECT  2.395 1.480 2.945 1.650 ;
        RECT  1.710 1.040 2.840 1.225 ;
        RECT  2.225 1.480 2.395 1.910 ;
        RECT  1.695 0.660 1.710 1.225 ;
        RECT  1.525 0.660 1.695 1.985 ;
        RECT  1.215 0.420 1.355 1.590 ;
        RECT  0.975 0.800 1.215 0.940 ;
        RECT  0.975 1.450 1.215 1.590 ;
        RECT  0.805 0.460 0.975 0.940 ;
        RECT  0.805 1.450 0.975 1.920 ;
        RECT  0.255 0.800 0.805 0.940 ;
        RECT  0.255 1.450 0.805 1.590 ;
        RECT  0.085 0.465 0.255 0.940 ;
        RECT  0.085 1.450 0.255 1.920 ;
    END
END ADDFHX4AD
MACRO ADDFHXLAD
    CLASS CORE ;
    FOREIGN ADDFHXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.350 0.735 7.490 1.675 ;
        RECT  7.305 0.735 7.350 0.905 ;
        RECT  7.305 1.505 7.350 1.675 ;
        END
        AntennaDiffArea 0.138 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.770 1.145 6.930 1.660 ;
        RECT  6.595 0.740 6.770 1.660 ;
        END
        AntennaDiffArea 0.151 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.265 0.970 6.445 1.380 ;
        RECT  6.215 1.140 6.265 1.380 ;
        END
        AntennaGateArea 0.0698 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.380 0.915 3.570 1.400 ;
        END
        AntennaGateArea 0.2574 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.050 0.440 1.310 ;
        RECT  0.070 0.905 0.210 1.375 ;
        END
        AntennaGateArea 0.1263 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.095 -0.210 7.560 0.210 ;
        RECT  6.925 -0.210 7.095 0.465 ;
        RECT  6.225 -0.210 6.925 0.210 ;
        RECT  5.965 -0.210 6.225 0.320 ;
        RECT  4.015 -0.210 5.965 0.210 ;
        RECT  3.755 -0.210 4.015 0.300 ;
        RECT  1.050 -0.210 3.755 0.210 ;
        RECT  0.530 -0.210 1.050 0.300 ;
        RECT  0.000 -0.210 0.530 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.120 2.310 7.560 2.730 ;
        RECT  6.950 2.075 7.120 2.730 ;
        RECT  6.025 2.310 6.950 2.730 ;
        RECT  5.765 2.220 6.025 2.730 ;
        RECT  3.615 2.310 5.765 2.730 ;
        RECT  3.355 2.020 3.615 2.730 ;
        RECT  0.950 2.310 3.355 2.730 ;
        RECT  0.950 1.965 1.010 2.135 ;
        RECT  0.650 1.965 0.950 2.730 ;
        RECT  0.580 1.965 0.650 2.135 ;
        RECT  0.000 2.310 0.650 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  7.170 1.020 7.230 1.280 ;
        RECT  7.050 1.020 7.170 1.900 ;
        RECT  6.505 1.780 7.050 1.900 ;
        RECT  6.295 2.020 6.830 2.140 ;
        RECT  6.390 0.390 6.560 0.560 ;
        RECT  6.385 1.740 6.505 1.900 ;
        RECT  6.095 1.500 6.435 1.620 ;
        RECT  6.145 0.440 6.390 0.560 ;
        RECT  5.125 1.740 6.385 1.860 ;
        RECT  6.175 1.980 6.295 2.140 ;
        RECT  5.555 1.980 6.175 2.100 ;
        RECT  6.095 0.440 6.145 1.030 ;
        RECT  6.025 0.440 6.095 1.620 ;
        RECT  5.075 0.440 6.025 0.560 ;
        RECT  5.975 0.910 6.025 1.620 ;
        RECT  5.675 1.180 5.975 1.350 ;
        RECT  5.765 0.680 5.905 0.800 ;
        RECT  5.645 0.680 5.765 1.060 ;
        RECT  5.555 0.940 5.645 1.060 ;
        RECT  5.555 1.500 5.645 1.620 ;
        RECT  5.435 0.940 5.555 1.620 ;
        RECT  5.465 1.980 5.555 2.140 ;
        RECT  5.315 0.700 5.525 0.820 ;
        RECT  4.595 2.020 5.465 2.140 ;
        RECT  5.385 1.500 5.435 1.620 ;
        RECT  5.195 0.700 5.315 1.355 ;
        RECT  5.125 1.235 5.195 1.355 ;
        RECT  5.005 1.235 5.125 1.860 ;
        RECT  4.955 0.440 5.075 1.115 ;
        RECT  4.835 0.995 4.955 1.115 ;
        RECT  4.715 0.375 4.835 0.635 ;
        RECT  4.715 0.995 4.835 1.875 ;
        RECT  4.595 0.755 4.785 0.875 ;
        RECT  4.115 0.420 4.715 0.555 ;
        RECT  4.475 0.755 4.595 2.140 ;
        RECT  4.075 2.020 4.475 2.140 ;
        RECT  4.235 0.685 4.355 1.900 ;
        RECT  3.930 1.780 4.235 1.900 ;
        RECT  3.995 0.420 4.115 1.660 ;
        RECT  3.655 0.420 3.995 0.555 ;
        RECT  3.760 1.780 3.930 2.095 ;
        RECT  3.755 0.675 3.875 1.300 ;
        RECT  3.355 1.780 3.760 1.900 ;
        RECT  3.445 0.675 3.755 0.795 ;
        RECT  3.550 0.380 3.655 0.555 ;
        RECT  2.570 0.380 3.550 0.500 ;
        RECT  3.330 0.620 3.445 0.795 ;
        RECT  3.235 1.640 3.355 1.900 ;
        RECT  2.810 0.620 3.330 0.740 ;
        RECT  3.115 0.860 3.225 0.980 ;
        RECT  2.995 0.860 3.115 2.140 ;
        RECT  2.965 0.860 2.995 0.980 ;
        RECT  1.535 2.020 2.995 2.140 ;
        RECT  2.810 1.170 2.875 1.900 ;
        RECT  2.755 0.620 2.810 1.900 ;
        RECT  2.690 0.620 2.755 1.290 ;
        RECT  1.915 1.780 2.755 1.900 ;
        RECT  2.570 1.400 2.635 1.660 ;
        RECT  2.450 0.380 2.570 1.660 ;
        RECT  2.210 0.385 2.330 1.650 ;
        RECT  1.600 0.385 2.210 0.505 ;
        RECT  2.130 1.480 2.210 1.650 ;
        RECT  1.915 0.660 1.995 0.830 ;
        RECT  1.795 0.660 1.915 1.900 ;
        RECT  1.535 0.660 1.635 0.830 ;
        RECT  1.480 0.385 1.600 0.540 ;
        RECT  1.415 0.660 1.535 2.140 ;
        RECT  0.680 0.420 1.480 0.540 ;
        RECT  1.175 1.130 1.295 1.680 ;
        RECT  0.975 1.430 1.175 1.680 ;
        RECT  0.800 0.770 0.975 1.680 ;
        RECT  0.560 0.420 0.680 1.615 ;
        RECT  0.085 0.615 0.560 0.785 ;
        RECT  0.230 1.495 0.560 1.615 ;
        RECT  0.110 1.495 0.230 1.790 ;
    END
END ADDFHXLAD
MACRO ADDFX1AD
    CLASS CORE ;
    FOREIGN ADDFX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.385 0.615 6.415 0.785 ;
        RECT  6.265 0.615 6.385 1.795 ;
        RECT  5.910 0.615 6.265 0.785 ;
        RECT  6.030 1.625 6.265 1.795 ;
        END
        AntennaDiffArea 0.2 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.790 0.575 6.930 1.920 ;
        RECT  6.745 0.575 6.790 0.745 ;
        RECT  6.770 1.400 6.790 1.920 ;
        END
        AntennaDiffArea 0.207 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.170 1.190 4.565 1.380 ;
        END
        AntennaGateArea 0.1093 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.205 1.055 0.490 1.375 ;
        RECT  0.070 1.145 0.205 1.375 ;
        END
        AntennaGateArea 0.14 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.985 0.910 2.505 1.130 ;
        END
        AntennaGateArea 0.1404 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.580 -0.210 7.000 0.210 ;
        RECT  6.320 -0.210 6.580 0.495 ;
        RECT  4.845 -0.210 6.320 0.210 ;
        RECT  4.585 -0.210 4.845 0.310 ;
        RECT  2.305 -0.210 4.585 0.210 ;
        RECT  2.185 -0.210 2.305 0.550 ;
        RECT  0.615 -0.210 2.185 0.210 ;
        RECT  0.445 -0.210 0.615 0.615 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.580 2.310 7.000 2.730 ;
        RECT  6.320 2.220 6.580 2.730 ;
        RECT  4.625 2.310 6.320 2.730 ;
        RECT  4.455 2.070 4.625 2.730 ;
        RECT  2.475 2.310 4.455 2.730 ;
        RECT  2.215 2.220 2.475 2.730 ;
        RECT  0.615 2.310 2.215 2.730 ;
        RECT  0.445 1.985 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.630 0.950 6.670 1.210 ;
        RECT  6.510 0.950 6.630 2.070 ;
        RECT  6.145 1.950 6.510 2.070 ;
        RECT  6.025 0.905 6.145 1.505 ;
        RECT  6.025 1.950 6.145 2.140 ;
        RECT  5.780 0.905 6.025 1.025 ;
        RECT  5.860 1.385 6.025 1.505 ;
        RECT  4.875 2.020 6.025 2.140 ;
        RECT  5.505 1.145 5.905 1.265 ;
        RECT  5.740 1.385 5.860 1.900 ;
        RECT  5.660 0.390 5.780 1.025 ;
        RECT  5.690 1.730 5.740 1.900 ;
        RECT  5.130 0.390 5.660 0.510 ;
        RECT  5.505 1.765 5.545 1.885 ;
        RECT  5.385 0.630 5.505 1.885 ;
        RECT  5.230 0.630 5.385 0.750 ;
        RECT  5.285 1.765 5.385 1.885 ;
        RECT  5.010 0.390 5.130 0.550 ;
        RECT  5.095 1.260 5.115 1.900 ;
        RECT  4.995 0.670 5.095 1.900 ;
        RECT  4.480 0.430 5.010 0.550 ;
        RECT  4.975 0.670 4.995 1.380 ;
        RECT  4.260 0.670 4.975 0.790 ;
        RECT  4.755 1.830 4.875 2.140 ;
        RECT  4.710 0.950 4.830 1.665 ;
        RECT  3.955 1.830 4.755 1.950 ;
        RECT  4.445 0.950 4.710 1.070 ;
        RECT  4.245 1.540 4.710 1.665 ;
        RECT  4.360 0.380 4.480 0.550 ;
        RECT  4.185 0.925 4.445 1.070 ;
        RECT  3.145 0.380 4.360 0.500 ;
        RECT  4.140 0.620 4.260 0.790 ;
        RECT  4.075 1.540 4.245 1.710 ;
        RECT  3.390 0.620 4.140 0.740 ;
        RECT  3.955 0.895 4.040 1.065 ;
        RECT  3.835 0.895 3.955 2.140 ;
        RECT  3.565 2.020 3.835 2.140 ;
        RECT  3.595 0.890 3.715 1.900 ;
        RECT  3.510 0.890 3.595 1.060 ;
        RECT  3.420 1.780 3.595 1.900 ;
        RECT  3.390 1.240 3.475 1.500 ;
        RECT  3.250 1.780 3.420 2.100 ;
        RECT  3.270 0.620 3.390 1.660 ;
        RECT  3.040 1.540 3.270 1.660 ;
        RECT  1.785 1.980 3.250 2.100 ;
        RECT  2.785 1.160 3.150 1.420 ;
        RECT  3.025 0.380 3.145 0.890 ;
        RECT  3.035 1.540 3.040 1.715 ;
        RECT  2.870 1.540 3.035 1.860 ;
        RECT  2.545 0.380 3.025 0.500 ;
        RECT  1.785 1.740 2.870 1.860 ;
        RECT  2.725 0.620 2.785 1.420 ;
        RECT  2.665 0.620 2.725 1.620 ;
        RECT  2.465 1.250 2.665 1.620 ;
        RECT  2.425 0.380 2.545 0.790 ;
        RECT  2.025 1.250 2.465 1.370 ;
        RECT  2.065 0.670 2.425 0.790 ;
        RECT  1.945 0.380 2.065 0.790 ;
        RECT  1.905 1.250 2.025 1.600 ;
        RECT  1.210 0.380 1.945 0.500 ;
        RECT  1.825 1.250 1.905 1.370 ;
        RECT  1.705 0.625 1.825 1.370 ;
        RECT  1.665 1.490 1.785 1.860 ;
        RECT  1.665 1.980 1.785 2.140 ;
        RECT  1.690 0.625 1.705 0.885 ;
        RECT  1.575 1.490 1.665 1.610 ;
        RECT  0.855 2.020 1.665 2.140 ;
        RECT  1.455 0.920 1.575 1.610 ;
        RECT  1.095 1.730 1.545 1.900 ;
        RECT  1.450 0.920 1.455 1.040 ;
        RECT  1.330 0.620 1.450 1.040 ;
        RECT  1.215 1.160 1.335 1.610 ;
        RECT  1.210 1.160 1.215 1.280 ;
        RECT  1.090 0.380 1.210 1.280 ;
        RECT  0.975 1.500 1.095 1.900 ;
        RECT  0.970 1.500 0.975 1.620 ;
        RECT  0.850 0.635 0.970 1.620 ;
        RECT  0.735 1.740 0.855 2.140 ;
        RECT  0.730 1.740 0.735 1.865 ;
        RECT  0.610 0.735 0.730 1.865 ;
        RECT  0.255 0.735 0.610 0.855 ;
        RECT  0.255 1.740 0.610 1.865 ;
        RECT  0.085 0.415 0.255 0.855 ;
        RECT  0.085 1.555 0.255 1.985 ;
    END
END ADDFX1AD
MACRO ADDFX2AD
    CLASS CORE ;
    FOREIGN ADDFX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.385 0.630 6.415 0.770 ;
        RECT  6.265 0.630 6.385 1.755 ;
        RECT  6.155 0.630 6.265 0.770 ;
        RECT  5.980 1.635 6.265 1.755 ;
        RECT  5.985 0.340 6.155 0.770 ;
        END
        AntennaDiffArea 0.373 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.790 0.330 6.930 2.190 ;
        RECT  6.760 0.330 6.790 0.850 ;
        RECT  6.760 1.410 6.790 2.190 ;
        END
        AntennaDiffArea 0.373 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.170 1.190 4.565 1.380 ;
        END
        AntennaGateArea 0.126 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.205 1.055 0.490 1.375 ;
        RECT  0.070 1.145 0.205 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.985 0.910 2.505 1.130 ;
        END
        AntennaGateArea 0.163 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.535 -0.210 7.000 0.210 ;
        RECT  6.365 -0.210 6.535 0.495 ;
        RECT  4.845 -0.210 6.365 0.210 ;
        RECT  4.585 -0.210 4.845 0.260 ;
        RECT  2.305 -0.210 4.585 0.210 ;
        RECT  2.185 -0.210 2.305 0.550 ;
        RECT  0.615 -0.210 2.185 0.210 ;
        RECT  0.445 -0.210 0.615 0.615 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.600 2.310 7.000 2.730 ;
        RECT  6.340 2.115 6.600 2.730 ;
        RECT  4.625 2.310 6.340 2.730 ;
        RECT  4.455 2.070 4.625 2.730 ;
        RECT  2.475 2.310 4.455 2.730 ;
        RECT  2.215 2.220 2.475 2.730 ;
        RECT  0.615 2.310 2.215 2.730 ;
        RECT  0.445 1.985 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.630 1.005 6.670 1.265 ;
        RECT  6.510 1.005 6.630 1.995 ;
        RECT  6.100 1.875 6.510 1.995 ;
        RECT  6.025 0.905 6.145 1.515 ;
        RECT  5.980 1.875 6.100 2.140 ;
        RECT  5.790 0.905 6.025 1.025 ;
        RECT  5.855 1.395 6.025 1.515 ;
        RECT  4.865 2.020 5.980 2.140 ;
        RECT  5.505 1.155 5.905 1.275 ;
        RECT  5.735 1.395 5.855 1.900 ;
        RECT  5.670 0.380 5.790 1.025 ;
        RECT  5.685 1.730 5.735 1.900 ;
        RECT  3.145 0.380 5.670 0.500 ;
        RECT  5.385 0.630 5.505 1.900 ;
        RECT  5.235 0.630 5.385 0.750 ;
        RECT  5.325 1.730 5.385 1.900 ;
        RECT  4.990 0.620 5.110 1.900 ;
        RECT  3.390 0.620 4.990 0.740 ;
        RECT  4.745 1.830 4.865 2.140 ;
        RECT  4.710 0.925 4.830 1.665 ;
        RECT  3.955 1.830 4.745 1.950 ;
        RECT  4.185 0.925 4.710 1.045 ;
        RECT  4.245 1.540 4.710 1.665 ;
        RECT  4.075 1.540 4.245 1.710 ;
        RECT  3.955 0.895 4.040 1.065 ;
        RECT  3.835 0.895 3.955 2.140 ;
        RECT  3.565 2.020 3.835 2.140 ;
        RECT  3.595 0.890 3.715 1.900 ;
        RECT  3.510 0.890 3.595 1.060 ;
        RECT  3.420 1.780 3.595 1.900 ;
        RECT  3.390 1.240 3.475 1.500 ;
        RECT  3.250 1.780 3.420 2.100 ;
        RECT  3.270 0.620 3.390 1.660 ;
        RECT  3.040 1.540 3.270 1.660 ;
        RECT  1.785 1.980 3.250 2.100 ;
        RECT  2.785 1.160 3.150 1.420 ;
        RECT  3.025 0.380 3.145 0.890 ;
        RECT  2.870 1.540 3.040 1.860 ;
        RECT  2.545 0.380 3.025 0.500 ;
        RECT  1.785 1.740 2.870 1.860 ;
        RECT  2.725 0.620 2.785 1.420 ;
        RECT  2.665 0.620 2.725 1.620 ;
        RECT  2.465 1.250 2.665 1.620 ;
        RECT  2.425 0.380 2.545 0.790 ;
        RECT  2.025 1.250 2.465 1.370 ;
        RECT  2.065 0.670 2.425 0.790 ;
        RECT  1.945 0.380 2.065 0.790 ;
        RECT  1.905 1.250 2.025 1.600 ;
        RECT  1.210 0.380 1.945 0.500 ;
        RECT  1.825 1.250 1.905 1.370 ;
        RECT  1.705 0.625 1.825 1.370 ;
        RECT  1.665 1.490 1.785 1.860 ;
        RECT  1.665 1.980 1.785 2.140 ;
        RECT  1.575 1.490 1.665 1.610 ;
        RECT  0.855 2.020 1.665 2.140 ;
        RECT  1.455 0.920 1.575 1.610 ;
        RECT  1.095 1.730 1.545 1.900 ;
        RECT  1.450 0.920 1.455 1.040 ;
        RECT  1.330 0.620 1.450 1.040 ;
        RECT  1.215 1.160 1.335 1.610 ;
        RECT  1.210 1.160 1.215 1.280 ;
        RECT  1.090 0.380 1.210 1.280 ;
        RECT  0.975 1.500 1.095 1.900 ;
        RECT  0.970 1.500 0.975 1.620 ;
        RECT  0.850 0.635 0.970 1.620 ;
        RECT  0.735 1.740 0.855 2.140 ;
        RECT  0.730 1.740 0.735 1.865 ;
        RECT  0.610 0.735 0.730 1.865 ;
        RECT  0.255 0.735 0.610 0.855 ;
        RECT  0.255 1.740 0.610 1.865 ;
        RECT  0.085 0.360 0.255 0.855 ;
        RECT  0.085 1.495 0.255 2.185 ;
    END
END ADDFX2AD
MACRO ADDFX4AD
    CLASS CORE ;
    FOREIGN ADDFX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.500 0.355 6.670 1.580 ;
        END
        AntennaDiffArea 0.422 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.390 0.725 7.490 1.515 ;
        RECT  7.350 0.355 7.390 2.170 ;
        RECT  7.220 0.355 7.350 0.895 ;
        RECT  7.220 1.345 7.350 2.170 ;
        END
        AntennaDiffArea 0.422 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.225 1.190 4.735 1.385 ;
        END
        AntennaGateArea 0.1268 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.045 0.420 1.215 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.980 0.910 2.500 1.130 ;
        END
        AntennaGateArea 0.1634 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.750 -0.210 7.840 0.210 ;
        RECT  7.580 -0.210 7.750 0.605 ;
        RECT  7.030 -0.210 7.580 0.210 ;
        RECT  6.860 -0.210 7.030 0.785 ;
        RECT  6.310 -0.210 6.860 0.210 ;
        RECT  6.140 -0.210 6.310 0.785 ;
        RECT  4.980 -0.210 6.140 0.210 ;
        RECT  4.720 -0.210 4.980 0.350 ;
        RECT  2.300 -0.210 4.720 0.210 ;
        RECT  2.180 -0.210 2.300 0.550 ;
        RECT  0.615 -0.210 2.180 0.210 ;
        RECT  0.445 -0.210 0.615 0.455 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.750 2.310 7.840 2.730 ;
        RECT  7.580 1.635 7.750 2.730 ;
        RECT  7.030 2.310 7.580 2.730 ;
        RECT  6.860 1.940 7.030 2.730 ;
        RECT  6.285 2.310 6.860 2.730 ;
        RECT  6.025 2.250 6.285 2.730 ;
        RECT  4.755 2.310 6.025 2.730 ;
        RECT  4.585 2.110 4.755 2.730 ;
        RECT  2.485 2.310 4.585 2.730 ;
        RECT  2.225 2.260 2.485 2.730 ;
        RECT  0.615 2.310 2.225 2.730 ;
        RECT  0.445 1.985 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.840 2.520 ;
        LAYER M1 ;
        RECT  7.090 1.080 7.230 1.200 ;
        RECT  6.970 1.080 7.090 1.820 ;
        RECT  6.220 1.700 6.970 1.820 ;
        RECT  6.260 0.915 6.380 1.515 ;
        RECT  5.945 0.915 6.260 1.035 ;
        RECT  5.980 1.395 6.260 1.515 ;
        RECT  6.100 1.700 6.220 2.130 ;
        RECT  5.665 1.155 6.140 1.275 ;
        RECT  4.995 2.010 6.100 2.130 ;
        RECT  5.860 1.395 5.980 1.890 ;
        RECT  5.825 0.470 5.945 1.035 ;
        RECT  5.810 1.720 5.860 1.890 ;
        RECT  4.600 0.470 5.825 0.590 ;
        RECT  5.545 0.730 5.665 1.890 ;
        RECT  5.365 0.730 5.545 0.850 ;
        RECT  5.405 1.770 5.545 1.890 ;
        RECT  5.115 0.710 5.235 1.890 ;
        RECT  4.360 0.710 5.115 0.830 ;
        RECT  4.875 1.870 4.995 2.130 ;
        RECT  4.855 0.950 4.975 1.700 ;
        RECT  4.045 1.870 4.875 1.990 ;
        RECT  4.285 0.950 4.855 1.070 ;
        RECT  4.335 1.580 4.855 1.700 ;
        RECT  4.480 0.380 4.600 0.590 ;
        RECT  3.140 0.380 4.480 0.500 ;
        RECT  4.240 0.620 4.360 0.830 ;
        RECT  4.165 1.580 4.335 1.750 ;
        RECT  3.510 0.620 4.240 0.740 ;
        RECT  4.045 0.895 4.135 1.065 ;
        RECT  3.925 0.895 4.045 2.140 ;
        RECT  3.685 2.020 3.925 2.140 ;
        RECT  3.685 0.860 3.805 1.900 ;
        RECT  3.630 0.860 3.685 1.120 ;
        RECT  3.500 1.780 3.685 1.900 ;
        RECT  3.510 1.240 3.565 1.500 ;
        RECT  3.390 0.620 3.510 1.660 ;
        RECT  3.330 1.780 3.500 2.140 ;
        RECT  3.115 1.540 3.390 1.660 ;
        RECT  0.855 2.020 3.330 2.140 ;
        RECT  3.145 1.160 3.265 1.420 ;
        RECT  2.780 1.300 3.145 1.420 ;
        RECT  3.020 0.380 3.140 0.880 ;
        RECT  2.995 1.540 3.115 1.860 ;
        RECT  2.540 0.380 3.020 0.500 ;
        RECT  1.795 1.740 2.995 1.860 ;
        RECT  2.745 0.620 2.780 1.420 ;
        RECT  2.660 0.620 2.745 1.620 ;
        RECT  2.485 1.250 2.660 1.620 ;
        RECT  2.420 0.380 2.540 0.790 ;
        RECT  2.035 1.250 2.485 1.370 ;
        RECT  2.060 0.670 2.420 0.790 ;
        RECT  1.940 0.380 2.060 0.790 ;
        RECT  1.915 1.250 2.035 1.600 ;
        RECT  1.220 0.380 1.940 0.500 ;
        RECT  1.820 1.250 1.915 1.370 ;
        RECT  1.700 0.620 1.820 1.370 ;
        RECT  1.675 1.490 1.795 1.860 ;
        RECT  1.580 1.490 1.675 1.610 ;
        RECT  1.460 0.830 1.580 1.610 ;
        RECT  1.385 1.730 1.555 1.900 ;
        RECT  1.340 0.620 1.460 0.950 ;
        RECT  1.095 1.730 1.385 1.850 ;
        RECT  1.220 1.150 1.340 1.610 ;
        RECT  1.100 0.380 1.220 1.270 ;
        RECT  0.980 1.505 1.095 1.850 ;
        RECT  0.975 0.560 0.980 1.850 ;
        RECT  0.860 0.560 0.975 1.625 ;
        RECT  0.735 1.745 0.855 2.140 ;
        RECT  0.710 1.745 0.735 1.865 ;
        RECT  0.590 0.760 0.710 1.865 ;
        RECT  0.465 0.760 0.590 0.880 ;
        RECT  0.255 1.745 0.590 1.865 ;
        RECT  0.345 0.575 0.465 0.880 ;
        RECT  0.085 0.575 0.345 0.745 ;
        RECT  0.085 1.570 0.255 2.000 ;
    END
END ADDFX4AD
MACRO ADDFXLAD
    CLASS CORE ;
    FOREIGN ADDFXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.385 0.615 6.415 0.785 ;
        RECT  6.265 0.615 6.385 1.745 ;
        RECT  5.910 0.615 6.265 0.785 ;
        RECT  5.985 1.625 6.265 1.745 ;
        END
        AntennaDiffArea 0.138 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.790 0.615 6.930 1.670 ;
        RECT  6.745 0.615 6.790 0.785 ;
        RECT  6.745 1.500 6.790 1.670 ;
        END
        AntennaDiffArea 0.138 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.170 1.190 4.565 1.380 ;
        END
        AntennaGateArea 0.1093 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.205 1.055 0.490 1.375 ;
        RECT  0.070 1.145 0.205 1.375 ;
        END
        AntennaGateArea 0.14 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.985 0.910 2.505 1.130 ;
        END
        AntennaGateArea 0.1404 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.580 -0.210 7.000 0.210 ;
        RECT  6.320 -0.210 6.580 0.495 ;
        RECT  4.845 -0.210 6.320 0.210 ;
        RECT  4.585 -0.210 4.845 0.310 ;
        RECT  2.305 -0.210 4.585 0.210 ;
        RECT  2.185 -0.210 2.305 0.550 ;
        RECT  0.615 -0.210 2.185 0.210 ;
        RECT  0.445 -0.210 0.615 0.615 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.580 2.310 7.000 2.730 ;
        RECT  6.320 2.220 6.580 2.730 ;
        RECT  4.625 2.310 6.320 2.730 ;
        RECT  4.455 2.070 4.625 2.730 ;
        RECT  2.475 2.310 4.455 2.730 ;
        RECT  2.215 2.220 2.475 2.730 ;
        RECT  0.615 2.310 2.215 2.730 ;
        RECT  0.445 1.985 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.625 0.950 6.670 1.210 ;
        RECT  6.505 0.950 6.625 2.070 ;
        RECT  6.145 1.950 6.505 2.070 ;
        RECT  6.025 0.905 6.145 1.505 ;
        RECT  6.025 1.950 6.145 2.140 ;
        RECT  5.780 0.905 6.025 1.025 ;
        RECT  5.860 1.385 6.025 1.505 ;
        RECT  4.875 2.020 6.025 2.140 ;
        RECT  5.505 1.145 5.905 1.265 ;
        RECT  5.740 1.385 5.860 1.900 ;
        RECT  5.660 0.390 5.780 1.025 ;
        RECT  5.690 1.730 5.740 1.900 ;
        RECT  5.130 0.390 5.660 0.510 ;
        RECT  5.505 1.765 5.545 1.885 ;
        RECT  5.385 0.630 5.505 1.885 ;
        RECT  5.230 0.630 5.385 0.750 ;
        RECT  5.285 1.765 5.385 1.885 ;
        RECT  5.010 0.390 5.130 0.550 ;
        RECT  5.095 1.260 5.115 1.900 ;
        RECT  4.995 0.670 5.095 1.900 ;
        RECT  4.480 0.430 5.010 0.550 ;
        RECT  4.975 0.670 4.995 1.380 ;
        RECT  4.260 0.670 4.975 0.790 ;
        RECT  4.755 1.830 4.875 2.140 ;
        RECT  4.710 0.925 4.830 1.665 ;
        RECT  3.955 1.830 4.755 1.950 ;
        RECT  4.185 0.925 4.710 1.045 ;
        RECT  4.245 1.540 4.710 1.665 ;
        RECT  4.360 0.380 4.480 0.550 ;
        RECT  3.145 0.380 4.360 0.500 ;
        RECT  4.140 0.620 4.260 0.790 ;
        RECT  4.075 1.540 4.245 1.710 ;
        RECT  3.390 0.620 4.140 0.740 ;
        RECT  3.955 0.895 4.040 1.065 ;
        RECT  3.835 0.895 3.955 2.140 ;
        RECT  3.565 2.020 3.835 2.140 ;
        RECT  3.595 0.890 3.715 1.900 ;
        RECT  3.510 0.890 3.595 1.060 ;
        RECT  3.420 1.780 3.595 1.900 ;
        RECT  3.390 1.240 3.475 1.500 ;
        RECT  3.250 1.780 3.420 2.100 ;
        RECT  3.270 0.620 3.390 1.660 ;
        RECT  3.040 1.540 3.270 1.660 ;
        RECT  1.785 1.980 3.250 2.100 ;
        RECT  2.785 1.160 3.150 1.420 ;
        RECT  3.025 0.380 3.145 0.890 ;
        RECT  2.870 1.540 3.040 1.860 ;
        RECT  2.545 0.380 3.025 0.500 ;
        RECT  1.785 1.740 2.870 1.860 ;
        RECT  2.725 0.620 2.785 1.420 ;
        RECT  2.665 0.620 2.725 1.620 ;
        RECT  2.465 1.250 2.665 1.620 ;
        RECT  2.425 0.380 2.545 0.790 ;
        RECT  2.025 1.250 2.465 1.370 ;
        RECT  2.065 0.670 2.425 0.790 ;
        RECT  1.945 0.380 2.065 0.790 ;
        RECT  1.905 1.250 2.025 1.600 ;
        RECT  1.210 0.380 1.945 0.500 ;
        RECT  1.825 1.250 1.905 1.370 ;
        RECT  1.705 0.625 1.825 1.370 ;
        RECT  1.665 1.490 1.785 1.860 ;
        RECT  1.665 1.980 1.785 2.140 ;
        RECT  1.690 0.625 1.705 0.885 ;
        RECT  1.575 1.490 1.665 1.610 ;
        RECT  0.855 2.020 1.665 2.140 ;
        RECT  1.455 0.920 1.575 1.610 ;
        RECT  1.095 1.730 1.545 1.900 ;
        RECT  1.450 0.920 1.455 1.040 ;
        RECT  1.330 0.620 1.450 1.040 ;
        RECT  1.215 1.160 1.335 1.610 ;
        RECT  1.210 1.160 1.215 1.280 ;
        RECT  1.090 0.380 1.210 1.280 ;
        RECT  0.975 1.500 1.095 1.900 ;
        RECT  0.970 1.500 0.975 1.620 ;
        RECT  0.850 0.635 0.970 1.620 ;
        RECT  0.735 1.740 0.855 2.140 ;
        RECT  0.730 1.740 0.735 1.865 ;
        RECT  0.610 0.735 0.730 1.865 ;
        RECT  0.255 0.735 0.610 0.855 ;
        RECT  0.255 1.740 0.610 1.865 ;
        RECT  0.085 0.415 0.255 0.855 ;
        RECT  0.085 1.555 0.255 1.985 ;
    END
END ADDFXLAD
MACRO ADDHX1AD
    CLASS CORE ;
    FOREIGN ADDHX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.735 0.865 1.890 1.375 ;
        RECT  1.675 0.650 1.735 1.620 ;
        RECT  1.605 0.650 1.675 1.895 ;
        RECT  1.555 1.500 1.605 1.895 ;
        RECT  1.505 1.725 1.555 1.895 ;
        END
        AntennaDiffArea 0.166 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.970 0.645 4.130 1.945 ;
        END
        AntennaDiffArea 0.207 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.710 0.360 1.880 0.530 ;
        RECT  1.480 0.410 1.710 0.530 ;
        RECT  1.375 0.410 1.480 1.385 ;
        RECT  1.360 0.410 1.375 1.610 ;
        RECT  1.145 1.190 1.360 1.610 ;
        END
        AntennaGateArea 0.1482 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.335 1.050 3.560 1.170 ;
        RECT  2.825 0.910 3.335 1.170 ;
        RECT  2.780 1.050 2.825 1.170 ;
        END
        AntennaGateArea 0.1494 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.720 -0.210 4.200 0.210 ;
        RECT  2.940 -0.210 3.720 0.300 ;
        RECT  0.630 -0.210 2.940 0.210 ;
        RECT  0.370 -0.210 0.630 0.300 ;
        RECT  0.000 -0.210 0.370 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.735 2.310 4.200 2.730 ;
        RECT  3.565 1.945 3.735 2.730 ;
        RECT  3.045 2.310 3.565 2.730 ;
        RECT  2.875 1.935 3.045 2.730 ;
        RECT  2.550 2.310 2.875 2.730 ;
        RECT  2.550 1.935 2.635 2.105 ;
        RECT  2.290 1.935 2.550 2.730 ;
        RECT  2.205 1.935 2.290 2.105 ;
        RECT  0.690 2.310 2.290 2.730 ;
        RECT  0.430 2.220 0.690 2.730 ;
        RECT  0.000 2.310 0.430 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  3.800 1.000 3.850 1.260 ;
        RECT  3.680 1.000 3.800 1.410 ;
        RECT  2.760 1.290 3.680 1.410 ;
        RECT  3.330 0.665 3.470 0.785 ;
        RECT  3.210 1.530 3.470 1.815 ;
        RECT  3.210 0.435 3.330 0.785 ;
        RECT  2.200 0.435 3.210 0.555 ;
        RECT  2.150 1.695 3.210 1.815 ;
        RECT  2.610 1.290 2.760 1.540 ;
        RECT  2.490 0.730 2.610 1.540 ;
        RECT  2.290 0.730 2.490 0.900 ;
        RECT  2.150 0.360 2.200 0.555 ;
        RECT  2.030 0.360 2.150 1.815 ;
        RECT  2.010 1.695 2.030 1.815 ;
        RECT  1.890 1.695 2.010 2.140 ;
        RECT  0.940 2.020 1.890 2.140 ;
        RECT  1.100 1.740 1.360 1.900 ;
        RECT  0.980 0.350 1.240 0.540 ;
        RECT  1.000 0.950 1.240 1.070 ;
        RECT  0.710 1.740 1.100 1.860 ;
        RECT  0.950 0.665 1.000 1.070 ;
        RECT  0.950 1.450 1.000 1.620 ;
        RECT  0.710 0.420 0.980 0.540 ;
        RECT  0.830 0.665 0.950 1.620 ;
        RECT  0.820 1.980 0.940 2.140 ;
        RECT  0.470 1.980 0.820 2.100 ;
        RECT  0.590 0.420 0.710 1.860 ;
        RECT  0.230 0.775 0.590 0.895 ;
        RECT  0.350 1.050 0.470 2.100 ;
        RECT  0.320 1.050 0.350 1.310 ;
        RECT  0.200 0.635 0.230 0.895 ;
        RECT  0.200 1.480 0.230 2.000 ;
        RECT  0.080 0.635 0.200 2.000 ;
    END
END ADDHX1AD
MACRO ADDHX2AD
    CLASS CORE ;
    FOREIGN ADDHX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 0.630 2.240 1.610 ;
        RECT  1.870 0.630 2.120 0.750 ;
        RECT  1.680 1.470 2.120 1.610 ;
        RECT  1.700 0.490 1.870 0.750 ;
        RECT  1.530 1.470 1.680 1.845 ;
        END
        AntennaDiffArea 0.368 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.370 4.410 2.035 ;
        END
        AntennaDiffArea 0.373 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.935 0.900 2.000 1.160 ;
        RECT  1.705 0.900 1.935 1.330 ;
        RECT  1.145 1.185 1.705 1.330 ;
        END
        AntennaGateArea 0.2718 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 1.040 3.630 1.160 ;
        RECT  2.850 0.865 3.010 1.160 ;
        END
        AntennaGateArea 0.3022 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.950 -0.210 4.480 0.210 ;
        RECT  3.690 -0.210 3.950 0.630 ;
        RECT  3.085 -0.210 3.690 0.210 ;
        RECT  2.915 -0.210 3.085 0.305 ;
        RECT  0.740 -0.210 2.915 0.210 ;
        RECT  0.480 -0.210 0.740 0.300 ;
        RECT  0.000 -0.210 0.480 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.920 2.310 4.480 2.730 ;
        RECT  3.750 1.810 3.920 2.730 ;
        RECT  3.040 2.310 3.750 2.730 ;
        RECT  2.260 2.220 3.040 2.730 ;
        RECT  0.740 2.310 2.260 2.730 ;
        RECT  0.480 2.220 0.740 2.730 ;
        RECT  0.000 2.310 0.480 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
        LAYER M1 ;
        RECT  4.010 0.750 4.130 1.685 ;
        RECT  3.440 0.750 4.010 0.870 ;
        RECT  3.465 1.565 4.010 1.685 ;
        RECT  3.770 1.010 3.890 1.445 ;
        RECT  2.835 1.325 3.770 1.445 ;
        RECT  3.295 1.565 3.465 2.050 ;
        RECT  3.320 0.440 3.440 0.870 ;
        RECT  2.775 0.440 3.320 0.560 ;
        RECT  2.050 1.930 3.295 2.050 ;
        RECT  2.480 1.325 2.835 1.530 ;
        RECT  2.655 0.390 2.775 0.560 ;
        RECT  2.015 0.390 2.655 0.510 ;
        RECT  2.360 0.665 2.480 1.530 ;
        RECT  1.880 1.730 2.050 2.160 ;
        RECT  0.480 1.980 1.880 2.100 ;
        RECT  1.325 0.395 1.495 0.565 ;
        RECT  0.720 1.740 1.375 1.860 ;
        RECT  0.965 0.750 1.360 0.970 ;
        RECT  0.720 0.445 1.325 0.565 ;
        RECT  0.840 0.750 0.965 1.620 ;
        RECT  0.600 0.445 0.720 1.860 ;
        RECT  0.240 0.725 0.600 0.845 ;
        RECT  0.360 1.025 0.480 2.100 ;
        RECT  0.330 1.025 0.360 1.285 ;
        RECT  0.190 0.370 0.240 0.890 ;
        RECT  0.190 1.510 0.240 2.030 ;
        RECT  0.120 0.370 0.190 2.030 ;
        RECT  0.070 0.725 0.120 2.030 ;
    END
END ADDHX2AD
MACRO ADDHX4AD
    CLASS CORE ;
    FOREIGN ADDHX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.015 0.650 3.275 0.895 ;
        RECT  2.435 1.460 3.155 1.580 ;
        RECT  2.505 0.770 3.015 0.895 ;
        RECT  2.450 0.435 2.505 0.895 ;
        RECT  2.310 0.435 2.450 0.955 ;
        RECT  2.245 1.460 2.435 1.620 ;
        RECT  1.875 0.775 2.310 0.895 ;
        RECT  1.875 1.500 2.245 1.620 ;
        RECT  1.755 0.620 1.875 1.620 ;
        RECT  1.550 0.620 1.755 0.740 ;
        RECT  1.450 1.500 1.755 1.620 ;
        END
        AntennaDiffArea 0.982 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.915 0.380 6.090 2.025 ;
        RECT  5.850 0.380 5.915 0.900 ;
        RECT  5.850 1.505 5.915 2.025 ;
        END
        AntennaDiffArea 0.422 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.060 1.015 3.230 1.330 ;
        RECT  2.125 1.180 3.060 1.330 ;
        RECT  2.005 1.110 2.125 1.370 ;
        END
        AntennaGateArea 0.5388 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.175 1.050 4.985 1.190 ;
        RECT  3.945 0.910 4.175 1.190 ;
        END
        AntennaGateArea 0.5918 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.330 -0.210 6.440 0.210 ;
        RECT  6.210 -0.210 6.330 0.880 ;
        RECT  5.635 -0.210 6.210 0.210 ;
        RECT  5.465 -0.210 5.635 0.530 ;
        RECT  4.930 -0.210 5.465 0.210 ;
        RECT  4.760 -0.210 4.930 0.270 ;
        RECT  4.190 -0.210 4.760 0.210 ;
        RECT  4.020 -0.210 4.190 0.550 ;
        RECT  1.040 -0.210 4.020 0.210 ;
        RECT  0.780 -0.210 1.040 0.260 ;
        RECT  0.255 -0.210 0.780 0.210 ;
        RECT  0.085 -0.210 0.255 0.845 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.330 2.310 6.440 2.730 ;
        RECT  6.210 1.510 6.330 2.730 ;
        RECT  5.635 2.310 6.210 2.730 ;
        RECT  5.465 1.895 5.635 2.730 ;
        RECT  4.950 2.310 5.465 2.730 ;
        RECT  4.780 1.795 4.950 2.730 ;
        RECT  4.210 2.310 4.780 2.730 ;
        RECT  4.040 2.200 4.210 2.730 ;
        RECT  3.400 2.310 4.040 2.730 ;
        RECT  3.230 1.985 3.400 2.730 ;
        RECT  0.995 2.310 3.230 2.730 ;
        RECT  0.825 2.265 0.995 2.730 ;
        RECT  0.255 2.310 0.825 2.730 ;
        RECT  0.085 1.890 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.440 2.520 ;
        LAYER M1 ;
        RECT  5.610 0.725 5.730 1.675 ;
        RECT  5.355 0.725 5.610 0.845 ;
        RECT  5.310 1.555 5.610 1.675 ;
        RECT  5.370 1.020 5.490 1.430 ;
        RECT  3.845 1.310 5.370 1.430 ;
        RECT  5.095 0.670 5.355 0.845 ;
        RECT  5.140 1.555 5.310 1.725 ;
        RECT  4.590 1.555 5.140 1.675 ;
        RECT  4.550 0.670 5.095 0.790 ;
        RECT  4.420 1.555 4.590 1.985 ;
        RECT  4.380 0.500 4.550 0.790 ;
        RECT  2.750 1.730 4.420 1.865 ;
        RECT  3.805 0.670 4.380 0.790 ;
        RECT  3.555 1.310 3.845 1.565 ;
        RECT  3.685 0.380 3.805 0.790 ;
        RECT  2.655 0.380 3.685 0.500 ;
        RECT  3.435 0.650 3.555 1.565 ;
        RECT  2.580 1.730 2.750 2.100 ;
        RECT  0.635 1.980 2.580 2.100 ;
        RECT  1.995 0.380 2.115 0.640 ;
        RECT  0.935 1.740 2.070 1.860 ;
        RECT  0.935 0.380 1.995 0.500 ;
        RECT  1.420 0.880 1.635 1.000 ;
        RECT  1.290 0.620 1.420 1.000 ;
        RECT  1.160 0.620 1.290 1.600 ;
        RECT  0.815 0.380 0.935 1.860 ;
        RECT  0.615 0.700 0.815 0.850 ;
        RECT  0.400 1.400 0.815 1.520 ;
        RECT  0.515 1.650 0.635 2.100 ;
        RECT  0.280 1.055 0.630 1.225 ;
        RECT  0.445 0.420 0.615 0.850 ;
        RECT  0.280 1.650 0.515 1.770 ;
        RECT  0.160 1.055 0.280 1.770 ;
    END
END ADDHX4AD
MACRO ADDHXLAD
    CLASS CORE ;
    FOREIGN ADDHXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.865 1.890 1.375 ;
        RECT  1.680 0.650 1.750 1.830 ;
        RECT  1.630 0.650 1.680 1.875 ;
        RECT  1.560 1.615 1.630 1.875 ;
        END
        AntennaDiffArea 0.112 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.990 0.735 4.130 1.680 ;
        RECT  3.935 0.735 3.990 0.905 ;
        RECT  3.960 1.420 3.990 1.680 ;
        END
        AntennaDiffArea 0.138 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.380 1.905 0.530 ;
        RECT  1.510 0.410 1.645 0.530 ;
        RECT  1.435 0.410 1.510 1.385 ;
        RECT  1.390 0.410 1.435 1.470 ;
        RECT  1.145 1.190 1.390 1.615 ;
        END
        AntennaGateArea 0.1315 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 0.865 3.290 1.165 ;
        RECT  2.750 1.045 2.870 1.165 ;
        END
        AntennaGateArea 0.1063 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.635 -0.210 4.200 0.210 ;
        RECT  3.115 -0.210 3.635 0.300 ;
        RECT  0.630 -0.210 3.115 0.210 ;
        RECT  0.370 -0.210 0.630 0.300 ;
        RECT  0.000 -0.210 0.370 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.725 2.310 4.200 2.730 ;
        RECT  3.555 1.875 3.725 2.730 ;
        RECT  3.035 2.310 3.555 2.730 ;
        RECT  2.865 1.910 3.035 2.730 ;
        RECT  2.415 2.310 2.865 2.730 ;
        RECT  2.245 1.910 2.415 2.730 ;
        RECT  0.690 2.310 2.245 2.730 ;
        RECT  0.430 2.220 0.690 2.730 ;
        RECT  0.000 2.310 0.430 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  3.800 1.065 3.865 1.235 ;
        RECT  3.680 1.065 3.800 1.440 ;
        RECT  2.725 1.320 3.680 1.440 ;
        RECT  3.340 0.625 3.480 0.745 ;
        RECT  3.415 1.585 3.460 1.705 ;
        RECT  3.200 1.585 3.415 1.790 ;
        RECT  3.220 0.435 3.340 0.745 ;
        RECT  2.195 0.435 3.220 0.555 ;
        RECT  2.145 1.670 3.200 1.790 ;
        RECT  2.610 1.320 2.725 1.550 ;
        RECT  2.490 0.735 2.610 1.550 ;
        RECT  2.305 0.735 2.490 0.905 ;
        RECT  2.145 0.360 2.195 0.555 ;
        RECT  2.040 0.360 2.145 1.790 ;
        RECT  2.025 0.360 2.040 2.140 ;
        RECT  1.920 1.615 2.025 2.140 ;
        RECT  0.935 2.020 1.920 2.140 ;
        RECT  1.100 1.740 1.360 1.900 ;
        RECT  1.010 0.345 1.270 0.540 ;
        RECT  1.000 0.945 1.240 1.065 ;
        RECT  0.710 1.740 1.100 1.860 ;
        RECT  0.710 0.420 1.010 0.540 ;
        RECT  0.950 0.660 1.000 1.065 ;
        RECT  0.950 1.450 1.000 1.620 ;
        RECT  0.830 0.660 0.950 1.620 ;
        RECT  0.815 1.980 0.935 2.140 ;
        RECT  0.470 1.980 0.815 2.100 ;
        RECT  0.590 0.420 0.710 1.860 ;
        RECT  0.280 0.830 0.590 0.950 ;
        RECT  0.350 1.070 0.470 2.100 ;
        RECT  0.230 0.690 0.280 0.950 ;
        RECT  0.110 0.690 0.230 1.770 ;
    END
END ADDHXLAD
MACRO AFCSHCINX2AD
    CLASS CORE ;
    FOREIGN AFCSHCINX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.850 0.790 15.890 1.540 ;
        RECT  15.750 0.365 15.850 2.030 ;
        RECT  15.730 0.365 15.750 0.940 ;
        RECT  15.730 1.390 15.750 2.030 ;
        END
        AntennaDiffArea 0.373 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  15.190 0.975 15.345 1.375 ;
        END
        AntennaGateArea 0.1762 ;
    END CS
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.220 0.620 10.335 0.880 ;
        RECT  10.220 1.145 10.290 1.375 ;
        RECT  10.100 0.620 10.220 2.015 ;
        END
        AntennaDiffArea 0.444 ;
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.890 0.860 9.005 0.980 ;
        RECT  8.835 0.860 8.890 1.095 ;
        RECT  8.715 0.860 8.835 1.900 ;
        END
        AntennaDiffArea 0.555 ;
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.275 1.190 13.055 1.385 ;
        END
        AntennaGateArea 0.3001 ;
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.135 1.080 6.395 1.250 ;
        RECT  5.920 1.080 6.135 1.375 ;
        RECT  5.705 1.080 5.920 1.250 ;
        END
        AntennaGateArea 0.2647 ;
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.195 0.865 4.410 1.255 ;
        END
        AntennaGateArea 0.4168 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.010 0.390 1.375 ;
        RECT  0.070 1.145 0.210 1.375 ;
        END
        AntennaGateArea 0.1605 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.515 -0.210 15.960 0.210 ;
        RECT  15.345 -0.210 15.515 0.700 ;
        RECT  14.805 -0.210 15.345 0.210 ;
        RECT  14.545 -0.210 14.805 0.565 ;
        RECT  13.535 -0.210 14.545 0.210 ;
        RECT  13.275 -0.210 13.535 0.300 ;
        RECT  12.180 -0.210 13.275 0.210 ;
        RECT  11.920 -0.210 12.180 0.300 ;
        RECT  6.915 -0.210 11.920 0.210 ;
        RECT  6.655 -0.210 6.915 0.415 ;
        RECT  6.165 -0.210 6.655 0.210 ;
        RECT  5.905 -0.210 6.165 0.380 ;
        RECT  4.545 -0.210 5.905 0.210 ;
        RECT  4.285 -0.210 4.545 0.300 ;
        RECT  1.330 -0.210 4.285 0.210 ;
        RECT  1.070 -0.210 1.330 0.300 ;
        RECT  0.680 -0.210 1.070 0.210 ;
        RECT  0.420 -0.210 0.680 0.300 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.560 2.310 15.960 2.730 ;
        RECT  15.300 2.130 15.560 2.730 ;
        RECT  14.895 2.310 15.300 2.730 ;
        RECT  14.635 2.030 14.895 2.730 ;
        RECT  13.405 2.310 14.635 2.730 ;
        RECT  12.885 2.230 13.405 2.730 ;
        RECT  12.275 2.310 12.885 2.730 ;
        RECT  12.015 2.220 12.275 2.730 ;
        RECT  5.735 2.310 12.015 2.730 ;
        RECT  5.475 2.105 5.735 2.730 ;
        RECT  4.725 2.310 5.475 2.730 ;
        RECT  4.465 2.220 4.725 2.730 ;
        RECT  1.260 2.310 4.465 2.730 ;
        RECT  1.140 2.195 1.260 2.730 ;
        RECT  0.615 2.310 1.140 2.730 ;
        RECT  0.445 1.735 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 15.960 2.520 ;
        LAYER M1 ;
        RECT  15.585 1.010 15.630 1.270 ;
        RECT  15.465 1.010 15.585 1.855 ;
        RECT  14.205 1.735 15.465 1.855 ;
        RECT  15.070 1.495 15.210 1.615 ;
        RECT  15.070 0.735 15.170 0.855 ;
        RECT  14.950 0.735 15.070 1.615 ;
        RECT  14.910 0.735 14.950 0.855 ;
        RECT  14.255 1.495 14.950 1.615 ;
        RECT  14.620 0.985 14.825 1.245 ;
        RECT  14.445 0.710 14.620 1.245 ;
        RECT  14.425 0.710 14.445 0.830 ;
        RECT  14.305 0.420 14.425 0.830 ;
        RECT  11.830 0.420 14.305 0.540 ;
        RECT  14.135 0.990 14.255 1.615 ;
        RECT  14.015 1.735 14.205 2.115 ;
        RECT  14.015 0.660 14.175 0.780 ;
        RECT  13.945 0.660 14.015 2.115 ;
        RECT  13.895 0.660 13.945 1.855 ;
        RECT  13.545 0.660 13.665 1.320 ;
        RECT  11.410 0.660 13.545 0.780 ;
        RECT  13.175 0.900 13.295 1.765 ;
        RECT  12.885 0.900 13.175 1.020 ;
        RECT  12.945 1.645 13.175 1.765 ;
        RECT  12.825 1.645 12.945 2.100 ;
        RECT  10.580 1.980 12.825 2.100 ;
        RECT  11.965 0.900 12.685 1.020 ;
        RECT  12.465 1.600 12.585 1.860 ;
        RECT  11.965 1.740 12.465 1.860 ;
        RECT  11.845 0.900 11.965 1.860 ;
        RECT  11.060 1.740 11.845 1.860 ;
        RECT  11.710 0.380 11.830 0.540 ;
        RECT  9.735 0.380 11.710 0.500 ;
        RECT  11.410 1.500 11.480 1.620 ;
        RECT  11.290 0.660 11.410 1.620 ;
        RECT  11.220 1.500 11.290 1.620 ;
        RECT  10.940 0.620 11.060 1.860 ;
        RECT  10.890 0.620 10.940 0.790 ;
        RECT  10.770 1.740 10.940 1.860 ;
        RECT  10.580 0.620 10.720 0.790 ;
        RECT  10.460 0.620 10.580 2.100 ;
        RECT  9.855 0.620 9.975 2.140 ;
        RECT  5.975 2.020 9.855 2.140 ;
        RECT  9.615 0.380 9.735 1.900 ;
        RECT  9.075 1.780 9.615 1.900 ;
        RECT  9.375 0.380 9.495 1.660 ;
        RECT  7.155 0.380 9.375 0.500 ;
        RECT  9.205 1.540 9.375 1.660 ;
        RECT  9.135 0.620 9.255 1.390 ;
        RECT  7.395 0.620 9.135 0.740 ;
        RECT  9.075 1.270 9.135 1.390 ;
        RECT  8.955 1.270 9.075 1.900 ;
        RECT  8.455 0.860 8.595 0.980 ;
        RECT  8.455 1.730 8.490 1.900 ;
        RECT  8.335 0.860 8.455 1.900 ;
        RECT  8.305 1.730 8.335 1.900 ;
        RECT  6.680 1.780 8.305 1.900 ;
        RECT  7.955 0.860 8.215 0.980 ;
        RECT  7.835 0.860 7.955 1.660 ;
        RECT  7.105 1.540 7.835 1.660 ;
        RECT  7.395 1.300 7.555 1.420 ;
        RECT  7.275 0.620 7.395 1.420 ;
        RECT  7.035 0.380 7.155 0.655 ;
        RECT  6.985 1.125 7.105 1.660 ;
        RECT  5.330 0.535 7.035 0.655 ;
        RECT  6.635 1.125 6.985 1.245 ;
        RECT  6.560 1.665 6.680 1.900 ;
        RECT  6.515 0.775 6.635 1.545 ;
        RECT  6.185 1.665 6.560 1.785 ;
        RECT  6.295 0.775 6.515 0.895 ;
        RECT  6.295 1.425 6.515 1.545 ;
        RECT  6.065 1.595 6.185 1.785 ;
        RECT  5.585 1.595 6.065 1.715 ;
        RECT  5.855 1.865 5.975 2.140 ;
        RECT  3.695 1.865 5.855 1.985 ;
        RECT  5.585 0.775 5.755 0.895 ;
        RECT  5.465 0.775 5.585 1.715 ;
        RECT  5.225 1.005 5.345 1.745 ;
        RECT  5.210 0.535 5.330 0.785 ;
        RECT  5.085 1.005 5.225 1.265 ;
        RECT  3.695 1.625 5.225 1.745 ;
        RECT  4.965 0.665 5.210 0.785 ;
        RECT  4.965 1.385 5.105 1.505 ;
        RECT  4.920 0.330 5.090 0.540 ;
        RECT  4.845 0.665 4.965 1.505 ;
        RECT  4.095 0.420 4.920 0.540 ;
        RECT  4.685 0.665 4.845 0.785 ;
        RECT  4.605 0.990 4.725 1.505 ;
        RECT  4.075 1.385 4.605 1.505 ;
        RECT  3.985 0.380 4.095 0.540 ;
        RECT  3.955 0.665 4.075 1.505 ;
        RECT  2.860 0.380 3.985 0.500 ;
        RECT  3.815 1.385 3.955 1.505 ;
        RECT  3.715 0.620 3.835 1.220 ;
        RECT  3.215 0.620 3.715 0.740 ;
        RECT  3.695 1.100 3.715 1.220 ;
        RECT  3.575 1.100 3.695 1.745 ;
        RECT  3.575 1.865 3.695 2.140 ;
        RECT  3.455 0.860 3.595 0.980 ;
        RECT  1.500 2.020 3.575 2.140 ;
        RECT  3.335 0.860 3.455 1.900 ;
        RECT  1.740 1.780 3.335 1.900 ;
        RECT  3.095 0.620 3.215 1.660 ;
        RECT  2.025 1.540 3.095 1.660 ;
        RECT  2.860 1.300 2.975 1.420 ;
        RECT  2.740 0.380 2.860 1.420 ;
        RECT  2.715 1.300 2.740 1.420 ;
        RECT  2.415 1.300 2.565 1.420 ;
        RECT  2.415 0.330 2.430 0.850 ;
        RECT  2.310 0.330 2.415 1.420 ;
        RECT  2.295 0.380 2.310 1.420 ;
        RECT  1.550 0.380 2.295 0.500 ;
        RECT  1.905 0.620 2.025 1.660 ;
        RECT  1.855 0.620 1.905 0.790 ;
        RECT  1.855 1.540 1.905 1.660 ;
        RECT  1.665 1.705 1.740 1.900 ;
        RECT  1.665 0.660 1.710 0.780 ;
        RECT  1.625 0.660 1.665 1.900 ;
        RECT  1.545 0.660 1.625 1.835 ;
        RECT  1.430 0.380 1.550 0.540 ;
        RECT  1.450 0.660 1.545 0.780 ;
        RECT  1.520 1.325 1.545 1.835 ;
        RECT  1.380 1.955 1.500 2.140 ;
        RECT  1.300 0.420 1.430 0.540 ;
        RECT  1.300 1.055 1.425 1.225 ;
        RECT  0.960 1.955 1.380 2.075 ;
        RECT  1.180 0.420 1.300 1.225 ;
        RECT  0.630 0.420 1.180 0.540 ;
        RECT  0.995 1.055 1.180 1.225 ;
        RECT  0.870 0.660 1.060 0.780 ;
        RECT  0.960 1.385 0.975 1.815 ;
        RECT  0.870 1.385 0.960 2.075 ;
        RECT  0.750 0.660 0.870 2.075 ;
        RECT  0.510 0.420 0.630 1.615 ;
        RECT  0.255 0.555 0.510 0.725 ;
        RECT  0.255 1.495 0.510 1.615 ;
        RECT  0.085 0.425 0.255 0.855 ;
        RECT  0.110 1.495 0.255 1.980 ;
        RECT  0.085 1.550 0.110 1.980 ;
    END
END AFCSHCINX2AD
MACRO AFCSHCINX4AD
    CLASS CORE ;
    FOREIGN AFCSHCINX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.410 0.790 16.450 1.540 ;
        RECT  16.310 0.365 16.410 2.030 ;
        RECT  16.290 0.365 16.310 0.940 ;
        RECT  16.290 1.390 16.310 2.030 ;
        END
        AntennaDiffArea 0.373 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  15.750 0.975 15.905 1.375 ;
        END
        AntennaGateArea 0.1761 ;
    END CS
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.850 0.620 10.895 0.880 ;
        RECT  10.780 0.620 10.850 1.690 ;
        RECT  10.710 0.620 10.780 2.015 ;
        RECT  10.660 1.495 10.710 2.015 ;
        END
        AntennaDiffArea 0.444 ;
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.405 0.860 9.565 0.980 ;
        RECT  9.285 0.860 9.405 1.900 ;
        RECT  9.275 1.285 9.285 1.900 ;
        RECT  9.030 1.285 9.275 1.795 ;
        END
        AntennaDiffArea 0.55 ;
    END CO0
    PIN CI1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  13.510 1.145 13.650 1.385 ;
        RECT  12.775 1.190 13.510 1.385 ;
        END
        AntennaGateArea 0.4267 ;
    END CI1N
    PIN CI0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.135 1.080 6.655 1.250 ;
        RECT  5.920 1.080 6.135 1.375 ;
        RECT  5.705 1.080 5.920 1.250 ;
        END
        AntennaGateArea 0.4265 ;
    END CI0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.195 0.865 4.410 1.255 ;
        END
        AntennaGateArea 0.4177 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.010 0.390 1.375 ;
        RECT  0.070 1.145 0.210 1.375 ;
        END
        AntennaGateArea 0.1605 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.075 -0.210 16.520 0.210 ;
        RECT  15.905 -0.210 16.075 0.700 ;
        RECT  15.480 -0.210 15.905 0.210 ;
        RECT  15.220 -0.210 15.480 0.500 ;
        RECT  14.220 -0.210 15.220 0.210 ;
        RECT  13.960 -0.210 14.220 0.300 ;
        RECT  13.460 -0.210 13.960 0.210 ;
        RECT  13.200 -0.210 13.460 0.300 ;
        RECT  12.730 -0.210 13.200 0.210 ;
        RECT  12.470 -0.210 12.730 0.300 ;
        RECT  7.505 -0.210 12.470 0.210 ;
        RECT  7.245 -0.210 7.505 0.380 ;
        RECT  6.805 -0.210 7.245 0.210 ;
        RECT  6.545 -0.210 6.805 0.380 ;
        RECT  6.085 -0.210 6.545 0.210 ;
        RECT  5.825 -0.210 6.085 0.380 ;
        RECT  4.545 -0.210 5.825 0.210 ;
        RECT  4.285 -0.210 4.545 0.300 ;
        RECT  1.330 -0.210 4.285 0.210 ;
        RECT  1.070 -0.210 1.330 0.300 ;
        RECT  0.680 -0.210 1.070 0.210 ;
        RECT  0.420 -0.210 0.680 0.300 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.120 2.310 16.520 2.730 ;
        RECT  15.860 2.130 16.120 2.730 ;
        RECT  15.480 2.310 15.860 2.730 ;
        RECT  15.220 2.030 15.480 2.730 ;
        RECT  14.120 2.310 15.220 2.730 ;
        RECT  13.950 1.960 14.120 2.730 ;
        RECT  13.425 2.310 13.950 2.730 ;
        RECT  13.165 2.230 13.425 2.730 ;
        RECT  12.775 2.310 13.165 2.730 ;
        RECT  12.515 2.220 12.775 2.730 ;
        RECT  5.480 2.310 12.515 2.730 ;
        RECT  5.220 2.140 5.480 2.730 ;
        RECT  4.625 2.310 5.220 2.730 ;
        RECT  4.455 2.150 4.625 2.730 ;
        RECT  1.260 2.310 4.455 2.730 ;
        RECT  1.140 2.195 1.260 2.730 ;
        RECT  0.615 2.310 1.140 2.730 ;
        RECT  0.445 1.735 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 16.520 2.520 ;
        LAYER M1 ;
        RECT  16.145 1.010 16.190 1.270 ;
        RECT  16.025 1.010 16.145 1.855 ;
        RECT  14.775 1.735 16.025 1.855 ;
        RECT  15.630 1.495 15.770 1.615 ;
        RECT  15.630 0.735 15.730 0.855 ;
        RECT  15.510 0.735 15.630 1.615 ;
        RECT  15.470 0.735 15.510 0.855 ;
        RECT  14.930 1.495 15.510 1.615 ;
        RECT  15.120 0.710 15.240 1.245 ;
        RECT  15.090 0.710 15.120 0.830 ;
        RECT  14.970 0.420 15.090 0.830 ;
        RECT  12.285 0.420 14.970 0.540 ;
        RECT  14.810 0.990 14.930 1.615 ;
        RECT  14.575 0.660 14.850 0.780 ;
        RECT  14.575 1.735 14.775 2.115 ;
        RECT  14.515 0.660 14.575 2.115 ;
        RECT  14.455 0.660 14.515 1.855 ;
        RECT  14.125 0.660 14.245 1.425 ;
        RECT  11.955 0.660 14.125 0.780 ;
        RECT  13.865 0.900 13.985 1.765 ;
        RECT  13.580 0.900 13.865 1.020 ;
        RECT  13.665 1.645 13.865 1.765 ;
        RECT  13.545 1.645 13.665 2.100 ;
        RECT  11.140 1.980 13.545 2.100 ;
        RECT  12.525 0.900 13.140 1.020 ;
        RECT  12.965 1.600 13.085 1.860 ;
        RECT  12.525 1.740 12.965 1.860 ;
        RECT  12.405 0.900 12.525 1.860 ;
        RECT  11.570 1.740 12.405 1.860 ;
        RECT  12.165 0.380 12.285 0.540 ;
        RECT  10.295 0.380 12.165 0.500 ;
        RECT  11.835 0.660 11.955 1.620 ;
        RECT  11.690 1.500 11.835 1.620 ;
        RECT  11.570 0.620 11.620 0.790 ;
        RECT  11.450 0.620 11.570 1.860 ;
        RECT  11.290 1.740 11.450 1.860 ;
        RECT  11.140 0.620 11.280 0.790 ;
        RECT  11.020 0.620 11.140 2.100 ;
        RECT  10.415 0.620 10.535 2.140 ;
        RECT  5.720 2.020 10.415 2.140 ;
        RECT  10.175 0.380 10.295 1.900 ;
        RECT  9.645 1.780 10.175 1.900 ;
        RECT  9.935 0.380 10.055 1.660 ;
        RECT  7.840 0.380 9.935 0.500 ;
        RECT  9.765 1.540 9.935 1.660 ;
        RECT  9.695 0.620 9.815 1.390 ;
        RECT  8.140 0.620 9.695 0.740 ;
        RECT  9.645 1.270 9.695 1.390 ;
        RECT  9.525 1.270 9.645 1.900 ;
        RECT  8.910 0.860 9.165 0.980 ;
        RECT  8.790 0.860 8.910 1.900 ;
        RECT  6.680 1.780 8.790 1.900 ;
        RECT  8.620 0.860 8.670 1.030 ;
        RECT  8.500 0.860 8.620 1.660 ;
        RECT  7.525 1.540 8.500 1.660 ;
        RECT  8.015 0.620 8.140 1.420 ;
        RECT  7.815 1.300 8.015 1.420 ;
        RECT  7.720 0.380 7.840 0.625 ;
        RECT  7.000 0.505 7.720 0.625 ;
        RECT  7.405 1.015 7.525 1.660 ;
        RECT  7.095 1.125 7.405 1.245 ;
        RECT  6.925 0.775 7.095 1.570 ;
        RECT  6.880 0.505 7.000 0.630 ;
        RECT  6.835 0.775 6.925 0.895 ;
        RECT  6.855 1.400 6.925 1.570 ;
        RECT  5.330 0.510 6.880 0.630 ;
        RECT  6.560 1.665 6.680 1.900 ;
        RECT  5.960 1.665 6.560 1.785 ;
        RECT  6.250 0.750 6.420 0.920 ;
        RECT  5.660 0.775 6.250 0.895 ;
        RECT  5.840 1.595 5.960 1.785 ;
        RECT  5.585 1.595 5.840 1.715 ;
        RECT  5.600 1.900 5.720 2.140 ;
        RECT  5.585 0.750 5.660 0.920 ;
        RECT  3.695 1.900 5.600 2.020 ;
        RECT  5.490 0.750 5.585 1.715 ;
        RECT  5.465 0.775 5.490 1.715 ;
        RECT  5.210 0.510 5.330 0.785 ;
        RECT  5.170 1.005 5.290 1.780 ;
        RECT  4.910 0.665 5.210 0.785 ;
        RECT  5.030 1.005 5.170 1.265 ;
        RECT  3.695 1.660 5.170 1.780 ;
        RECT  4.920 0.330 5.090 0.540 ;
        RECT  4.910 1.385 5.050 1.505 ;
        RECT  4.095 0.420 4.920 0.540 ;
        RECT  4.790 0.665 4.910 1.505 ;
        RECT  4.685 0.665 4.790 0.785 ;
        RECT  4.550 0.990 4.670 1.505 ;
        RECT  4.075 1.385 4.550 1.505 ;
        RECT  3.985 0.380 4.095 0.540 ;
        RECT  3.985 0.665 4.075 1.505 ;
        RECT  2.860 0.380 3.985 0.500 ;
        RECT  3.955 0.665 3.985 1.530 ;
        RECT  3.815 1.360 3.955 1.530 ;
        RECT  3.715 0.620 3.835 1.220 ;
        RECT  3.215 0.620 3.715 0.740 ;
        RECT  3.695 1.100 3.715 1.220 ;
        RECT  3.575 1.100 3.695 1.780 ;
        RECT  3.575 1.900 3.695 2.140 ;
        RECT  3.455 0.860 3.595 0.980 ;
        RECT  1.500 2.020 3.575 2.140 ;
        RECT  3.335 0.860 3.455 1.900 ;
        RECT  1.740 1.780 3.335 1.900 ;
        RECT  3.095 0.620 3.215 1.660 ;
        RECT  2.025 1.540 3.095 1.660 ;
        RECT  2.860 1.300 2.975 1.420 ;
        RECT  2.740 0.380 2.860 1.420 ;
        RECT  2.715 1.300 2.740 1.420 ;
        RECT  2.405 1.300 2.565 1.420 ;
        RECT  2.405 0.375 2.455 0.805 ;
        RECT  2.285 0.375 2.405 1.420 ;
        RECT  1.550 0.380 2.285 0.500 ;
        RECT  1.905 0.620 2.025 1.660 ;
        RECT  1.855 0.620 1.905 0.790 ;
        RECT  1.855 1.540 1.905 1.660 ;
        RECT  1.665 1.705 1.740 1.900 ;
        RECT  1.665 0.660 1.710 0.780 ;
        RECT  1.625 0.660 1.665 1.900 ;
        RECT  1.545 0.660 1.625 1.835 ;
        RECT  1.430 0.380 1.550 0.540 ;
        RECT  1.450 0.660 1.545 0.780 ;
        RECT  1.520 1.575 1.545 1.835 ;
        RECT  1.380 1.955 1.500 2.140 ;
        RECT  1.300 0.420 1.430 0.540 ;
        RECT  1.300 1.055 1.425 1.225 ;
        RECT  0.960 1.955 1.380 2.075 ;
        RECT  1.180 0.420 1.300 1.225 ;
        RECT  0.630 0.420 1.180 0.540 ;
        RECT  0.995 1.055 1.180 1.225 ;
        RECT  0.870 0.660 1.060 0.780 ;
        RECT  0.960 1.385 0.975 1.815 ;
        RECT  0.870 1.385 0.960 2.075 ;
        RECT  0.750 0.660 0.870 2.075 ;
        RECT  0.510 0.420 0.630 1.615 ;
        RECT  0.255 0.555 0.510 0.725 ;
        RECT  0.255 1.495 0.510 1.615 ;
        RECT  0.085 0.425 0.255 0.855 ;
        RECT  0.110 1.495 0.255 1.980 ;
        RECT  0.085 1.550 0.110 1.980 ;
    END
END AFCSHCINX4AD
MACRO AFCSHCONX2AD
    CLASS CORE ;
    FOREIGN AFCSHCONX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.035 0.730 15.050 1.685 ;
        RECT  14.910 0.440 15.035 1.975 ;
        RECT  14.865 0.440 14.910 0.870 ;
        RECT  14.865 1.545 14.910 1.975 ;
        END
        AntennaDiffArea 0.373 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.080 1.065 14.490 1.375 ;
        END
        AntennaGateArea 0.1764 ;
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.350 1.145 9.450 1.375 ;
        RECT  9.275 0.620 9.350 1.375 ;
        RECT  9.180 0.620 9.275 1.995 ;
        RECT  9.135 1.235 9.180 1.995 ;
        END
        AntennaDiffArea 0.451 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.865 0.860 7.975 0.980 ;
        RECT  7.745 0.860 7.865 1.900 ;
        RECT  7.695 0.860 7.745 1.655 ;
        RECT  7.630 1.145 7.695 1.655 ;
        END
        AntennaDiffArea 0.503 ;
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.495 1.160 12.015 1.380 ;
        END
        AntennaGateArea 0.3136 ;
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.070 4.980 1.375 ;
        END
        AntennaGateArea 0.2678 ;
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.055 0.360 1.225 ;
        RECT  0.070 1.055 0.210 1.375 ;
        END
        AntennaGateArea 0.4453 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 0.995 3.130 1.165 ;
        RECT  2.870 0.865 3.010 1.165 ;
        RECT  2.700 0.995 2.870 1.165 ;
        END
        AntennaGateArea 0.3179 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.675 -0.210 15.120 0.210 ;
        RECT  14.505 -0.210 14.675 0.870 ;
        RECT  13.880 -0.210 14.505 0.210 ;
        RECT  13.620 -0.210 13.880 0.630 ;
        RECT  12.555 -0.210 13.620 0.210 ;
        RECT  12.295 -0.210 12.555 0.260 ;
        RECT  11.345 -0.210 12.295 0.210 ;
        RECT  10.825 -0.210 11.345 0.260 ;
        RECT  6.015 -0.210 10.825 0.210 ;
        RECT  5.755 -0.210 6.015 0.415 ;
        RECT  5.220 -0.210 5.755 0.210 ;
        RECT  4.960 -0.210 5.220 0.415 ;
        RECT  2.965 -0.210 4.960 0.210 ;
        RECT  2.795 -0.210 2.965 0.720 ;
        RECT  1.290 -0.210 2.795 0.210 ;
        RECT  1.170 -0.210 1.290 0.840 ;
        RECT  0.660 -0.210 1.170 0.210 ;
        RECT  0.400 -0.210 0.660 0.670 ;
        RECT  0.000 -0.210 0.400 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.675 2.310 15.120 2.730 ;
        RECT  14.505 1.980 14.675 2.730 ;
        RECT  13.985 2.310 14.505 2.730 ;
        RECT  13.815 1.980 13.985 2.730 ;
        RECT  12.555 2.310 13.815 2.730 ;
        RECT  11.865 2.175 12.555 2.730 ;
        RECT  11.255 2.310 11.865 2.730 ;
        RECT  10.995 2.220 11.255 2.730 ;
        RECT  4.680 2.310 10.995 2.730 ;
        RECT  4.510 2.115 4.680 2.730 ;
        RECT  3.125 2.310 4.510 2.730 ;
        RECT  2.955 2.220 3.125 2.730 ;
        RECT  1.380 2.310 2.955 2.730 ;
        RECT  1.120 2.290 1.380 2.730 ;
        RECT  0.615 2.310 1.120 2.730 ;
        RECT  0.445 2.085 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 15.120 2.520 ;
        LAYER M1 ;
        RECT  14.625 1.020 14.745 1.860 ;
        RECT  13.225 1.740 14.625 1.860 ;
        RECT  14.080 0.740 14.340 0.870 ;
        RECT  13.960 1.500 14.340 1.620 ;
        RECT  13.960 0.750 14.080 0.870 ;
        RECT  13.840 0.750 13.960 1.620 ;
        RECT  13.340 1.385 13.840 1.505 ;
        RECT  13.580 1.035 13.720 1.155 ;
        RECT  13.475 0.780 13.580 1.155 ;
        RECT  13.460 0.380 13.475 1.155 ;
        RECT  13.355 0.380 13.460 0.900 ;
        RECT  8.725 0.380 13.355 0.500 ;
        RECT  13.220 1.020 13.340 1.505 ;
        RECT  13.055 1.655 13.225 2.085 ;
        RECT  13.080 1.020 13.220 1.140 ;
        RECT  12.955 0.660 13.175 0.830 ;
        RECT  12.955 1.655 13.055 1.860 ;
        RECT  12.835 0.660 12.955 1.860 ;
        RECT  12.595 0.620 12.715 1.380 ;
        RECT  10.410 0.620 12.595 0.740 ;
        RECT  12.135 0.860 12.255 1.945 ;
        RECT  11.915 0.860 12.135 0.980 ;
        RECT  11.295 1.825 12.135 1.945 ;
        RECT  11.375 0.860 11.795 0.980 ;
        RECT  11.375 1.585 11.635 1.705 ;
        RECT  11.255 0.860 11.375 1.705 ;
        RECT  11.175 1.825 11.295 2.100 ;
        RECT  10.955 1.585 11.255 1.705 ;
        RECT  9.710 1.980 11.175 2.100 ;
        RECT  10.885 1.065 10.955 1.705 ;
        RECT  10.835 1.065 10.885 1.860 ;
        RECT  10.765 1.585 10.835 1.860 ;
        RECT  10.000 1.740 10.765 1.860 ;
        RECT  10.410 1.500 10.555 1.620 ;
        RECT  10.290 0.620 10.410 1.620 ;
        RECT  10.240 0.660 10.290 0.830 ;
        RECT  10.000 0.620 10.050 0.790 ;
        RECT  9.880 0.620 10.000 1.860 ;
        RECT  9.590 0.620 9.710 2.100 ;
        RECT  9.540 0.620 9.590 0.790 ;
        RECT  9.470 1.520 9.590 2.100 ;
        RECT  8.965 1.085 9.015 2.140 ;
        RECT  8.895 0.620 8.965 2.140 ;
        RECT  8.845 0.620 8.895 1.205 ;
        RECT  4.950 2.020 8.895 2.140 ;
        RECT  8.725 1.315 8.775 1.900 ;
        RECT  8.655 0.380 8.725 1.900 ;
        RECT  8.605 0.380 8.655 1.435 ;
        RECT  8.105 1.780 8.655 1.900 ;
        RECT  8.485 1.535 8.515 1.655 ;
        RECT  8.365 0.380 8.485 1.655 ;
        RECT  6.275 0.380 8.365 0.500 ;
        RECT  8.255 1.535 8.365 1.655 ;
        RECT  8.125 0.620 8.245 1.410 ;
        RECT  6.545 0.620 8.125 0.740 ;
        RECT  8.105 1.290 8.125 1.410 ;
        RECT  7.985 1.290 8.105 1.900 ;
        RECT  7.435 0.860 7.575 0.980 ;
        RECT  7.435 1.730 7.530 1.900 ;
        RECT  7.315 0.860 7.435 1.900 ;
        RECT  5.700 1.780 7.315 1.900 ;
        RECT  7.055 0.860 7.195 0.980 ;
        RECT  6.935 0.860 7.055 1.660 ;
        RECT  5.985 1.540 6.935 1.660 ;
        RECT  6.425 0.620 6.545 1.420 ;
        RECT  6.275 1.300 6.425 1.420 ;
        RECT  6.155 0.380 6.275 0.655 ;
        RECT  4.410 0.535 6.155 0.655 ;
        RECT  5.650 1.005 5.985 1.265 ;
        RECT  5.865 1.435 5.985 1.660 ;
        RECT  5.650 1.435 5.865 1.555 ;
        RECT  5.580 1.675 5.700 1.900 ;
        RECT  5.390 0.780 5.650 1.555 ;
        RECT  5.185 1.675 5.580 1.795 ;
        RECT  5.305 1.435 5.390 1.555 ;
        RECT  5.065 1.525 5.185 1.795 ;
        RECT  4.430 1.525 5.065 1.645 ;
        RECT  4.830 1.840 4.950 2.140 ;
        RECT  4.430 0.775 4.840 0.895 ;
        RECT  4.285 1.840 4.830 1.960 ;
        RECT  4.310 0.775 4.430 1.645 ;
        RECT  4.290 0.380 4.410 0.655 ;
        RECT  3.480 0.380 4.290 0.500 ;
        RECT  4.165 1.840 4.285 2.100 ;
        RECT  2.440 1.980 4.165 2.100 ;
        RECT  3.930 0.620 4.050 1.745 ;
        RECT  3.840 1.040 3.930 1.300 ;
        RECT  3.600 0.620 3.720 1.860 ;
        RECT  3.010 1.740 3.600 1.860 ;
        RECT  3.360 0.380 3.480 1.620 ;
        RECT  3.155 0.380 3.360 0.810 ;
        RECT  2.890 1.590 3.010 1.860 ;
        RECT  2.340 1.590 2.890 1.710 ;
        RECT  2.580 1.350 2.770 1.470 ;
        RECT  2.460 0.380 2.580 1.470 ;
        RECT  1.610 0.380 2.460 0.500 ;
        RECT  2.320 1.830 2.440 2.100 ;
        RECT  2.220 0.630 2.340 1.710 ;
        RECT  2.020 1.830 2.320 1.950 ;
        RECT  1.820 0.630 2.220 0.750 ;
        RECT  2.130 1.590 2.220 1.710 ;
        RECT  1.800 2.070 2.200 2.190 ;
        RECT  1.980 1.120 2.100 1.470 ;
        RECT  1.900 1.760 2.020 1.950 ;
        RECT  1.385 1.350 1.980 1.470 ;
        RECT  0.600 1.760 1.900 1.880 ;
        RECT  1.680 2.020 1.800 2.190 ;
        RECT  1.210 2.020 1.680 2.140 ;
        RECT  1.490 0.380 1.610 1.210 ;
        RECT  1.080 1.090 1.490 1.210 ;
        RECT  1.265 1.350 1.385 1.540 ;
        RECT  1.020 1.420 1.265 1.540 ;
        RECT  0.950 2.020 1.210 2.150 ;
        RECT  0.960 1.015 1.080 1.275 ;
        RECT  0.840 1.420 1.020 1.620 ;
        RECT  0.840 0.390 0.975 0.895 ;
        RECT  0.805 0.390 0.840 1.620 ;
        RECT  0.760 0.775 0.805 1.620 ;
        RECT  0.720 0.775 0.760 1.540 ;
        RECT  0.480 0.790 0.600 1.880 ;
        RECT  0.255 0.790 0.480 0.910 ;
        RECT  0.255 1.760 0.480 1.880 ;
        RECT  0.085 0.395 0.255 0.910 ;
        RECT  0.085 1.595 0.255 2.025 ;
    END
END AFCSHCONX2AD
MACRO AFCSHCONX4AD
    CLASS CORE ;
    FOREIGN AFCSHCONX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.155 0.730 16.170 1.685 ;
        RECT  16.030 0.440 16.155 1.975 ;
        RECT  15.985 0.440 16.030 0.870 ;
        RECT  15.985 1.545 16.030 1.975 ;
        END
        AntennaDiffArea 0.373 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  15.365 0.990 15.610 1.375 ;
        END
        AntennaGateArea 0.1764 ;
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.470 1.005 10.570 1.515 ;
        RECT  10.395 0.620 10.470 1.515 ;
        RECT  10.300 0.620 10.395 1.995 ;
        RECT  10.255 1.235 10.300 1.995 ;
        END
        AntennaDiffArea 0.451 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.985 0.860 9.095 0.980 ;
        RECT  8.865 0.860 8.985 1.900 ;
        RECT  8.815 0.860 8.865 1.795 ;
        RECT  8.750 1.285 8.815 1.795 ;
        END
        AntennaDiffArea 0.503 ;
    END CO0N
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.615 1.160 13.135 1.380 ;
        END
        AntennaGateArea 0.5649 ;
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.540 1.095 5.890 1.215 ;
        RECT  5.110 1.070 5.540 1.375 ;
        END
        AntennaGateArea 0.6164 ;
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.055 0.360 1.225 ;
        RECT  0.070 1.055 0.210 1.375 ;
        END
        AntennaGateArea 0.4453 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 0.995 3.130 1.165 ;
        RECT  2.870 0.865 3.010 1.165 ;
        RECT  2.700 0.995 2.870 1.165 ;
        END
        AntennaGateArea 0.3179 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.795 -0.210 16.240 0.210 ;
        RECT  15.625 -0.210 15.795 0.870 ;
        RECT  15.000 -0.210 15.625 0.210 ;
        RECT  14.740 -0.210 15.000 0.630 ;
        RECT  13.630 -0.210 14.740 0.210 ;
        RECT  13.460 -0.210 13.630 0.255 ;
        RECT  12.995 -0.210 13.460 0.210 ;
        RECT  12.735 -0.210 12.995 0.260 ;
        RECT  12.205 -0.210 12.735 0.210 ;
        RECT  11.945 -0.210 12.205 0.260 ;
        RECT  7.135 -0.210 11.945 0.210 ;
        RECT  6.875 -0.210 7.135 0.415 ;
        RECT  6.345 -0.210 6.875 0.210 ;
        RECT  6.085 -0.210 6.345 0.415 ;
        RECT  5.260 -0.210 6.085 0.210 ;
        RECT  5.000 -0.210 5.260 0.415 ;
        RECT  4.500 -0.210 5.000 0.210 ;
        RECT  4.240 -0.210 4.500 0.415 ;
        RECT  2.965 -0.210 4.240 0.210 ;
        RECT  2.795 -0.210 2.965 0.720 ;
        RECT  1.290 -0.210 2.795 0.210 ;
        RECT  1.170 -0.210 1.290 0.840 ;
        RECT  0.660 -0.210 1.170 0.210 ;
        RECT  0.400 -0.210 0.660 0.670 ;
        RECT  0.000 -0.210 0.400 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.795 2.310 16.240 2.730 ;
        RECT  15.625 1.980 15.795 2.730 ;
        RECT  15.105 2.310 15.625 2.730 ;
        RECT  14.935 1.980 15.105 2.730 ;
        RECT  13.780 2.310 14.935 2.730 ;
        RECT  13.660 1.665 13.780 2.730 ;
        RECT  13.090 2.310 13.660 2.730 ;
        RECT  12.920 2.265 13.090 2.730 ;
        RECT  12.375 2.310 12.920 2.730 ;
        RECT  12.115 2.220 12.375 2.730 ;
        RECT  5.190 2.310 12.115 2.730 ;
        RECT  5.010 2.070 5.190 2.730 ;
        RECT  4.455 2.310 5.010 2.730 ;
        RECT  4.285 1.980 4.455 2.730 ;
        RECT  3.125 2.310 4.285 2.730 ;
        RECT  2.955 2.220 3.125 2.730 ;
        RECT  1.380 2.310 2.955 2.730 ;
        RECT  1.120 2.290 1.380 2.730 ;
        RECT  0.615 2.310 1.120 2.730 ;
        RECT  0.445 2.085 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 16.240 2.520 ;
        LAYER M1 ;
        RECT  15.745 1.020 15.865 1.860 ;
        RECT  14.415 1.740 15.745 1.860 ;
        RECT  15.245 0.740 15.460 0.870 ;
        RECT  15.245 1.500 15.460 1.620 ;
        RECT  15.200 0.740 15.245 1.620 ;
        RECT  15.125 0.750 15.200 1.620 ;
        RECT  14.460 1.385 15.125 1.505 ;
        RECT  14.730 0.780 14.850 1.240 ;
        RECT  14.595 0.780 14.730 0.900 ;
        RECT  14.475 0.380 14.595 0.900 ;
        RECT  9.845 0.380 14.475 0.500 ;
        RECT  14.340 1.020 14.460 1.505 ;
        RECT  14.245 1.655 14.415 2.085 ;
        RECT  14.200 1.020 14.340 1.140 ;
        RECT  14.075 0.660 14.295 0.830 ;
        RECT  14.075 1.655 14.245 1.860 ;
        RECT  13.955 0.660 14.075 1.860 ;
        RECT  13.715 0.620 13.835 1.380 ;
        RECT  11.530 0.620 13.715 0.740 ;
        RECT  13.255 0.860 13.375 2.100 ;
        RECT  13.115 0.860 13.255 0.980 ;
        RECT  10.830 1.980 13.255 2.100 ;
        RECT  12.475 1.585 12.755 1.705 ;
        RECT  12.475 0.860 12.615 0.980 ;
        RECT  12.355 0.860 12.475 1.705 ;
        RECT  12.075 1.585 12.355 1.705 ;
        RECT  12.005 1.065 12.075 1.705 ;
        RECT  11.955 1.065 12.005 1.860 ;
        RECT  11.885 1.585 11.955 1.860 ;
        RECT  11.120 1.740 11.885 1.860 ;
        RECT  11.530 1.500 11.675 1.620 ;
        RECT  11.410 0.620 11.530 1.620 ;
        RECT  11.360 0.660 11.410 0.830 ;
        RECT  11.120 0.620 11.170 0.790 ;
        RECT  11.000 0.620 11.120 1.860 ;
        RECT  10.710 0.620 10.830 2.100 ;
        RECT  10.660 0.620 10.710 0.790 ;
        RECT  10.590 1.690 10.710 2.100 ;
        RECT  10.085 1.085 10.135 2.140 ;
        RECT  10.015 0.620 10.085 2.140 ;
        RECT  9.965 0.620 10.015 1.205 ;
        RECT  5.430 2.020 10.015 2.140 ;
        RECT  9.845 1.315 9.895 1.900 ;
        RECT  9.775 0.380 9.845 1.900 ;
        RECT  9.725 0.380 9.775 1.435 ;
        RECT  9.225 1.780 9.775 1.900 ;
        RECT  9.605 1.535 9.635 1.655 ;
        RECT  9.485 0.380 9.605 1.655 ;
        RECT  7.395 0.380 9.485 0.500 ;
        RECT  9.375 1.535 9.485 1.655 ;
        RECT  9.245 0.620 9.365 1.410 ;
        RECT  7.665 0.620 9.245 0.740 ;
        RECT  9.225 1.290 9.245 1.410 ;
        RECT  9.105 1.290 9.225 1.900 ;
        RECT  8.555 0.860 8.695 0.980 ;
        RECT  8.555 1.640 8.625 1.900 ;
        RECT  8.435 0.860 8.555 1.900 ;
        RECT  6.540 1.780 8.435 1.900 ;
        RECT  8.175 0.860 8.315 0.980 ;
        RECT  8.055 0.860 8.175 1.660 ;
        RECT  7.105 1.540 8.055 1.660 ;
        RECT  7.545 0.620 7.665 1.420 ;
        RECT  7.395 1.300 7.545 1.420 ;
        RECT  7.275 0.380 7.395 0.655 ;
        RECT  3.990 0.535 7.275 0.655 ;
        RECT  6.985 1.005 7.105 1.660 ;
        RECT  6.440 1.075 6.985 1.195 ;
        RECT  6.440 0.780 6.725 0.900 ;
        RECT  6.405 1.435 6.650 1.555 ;
        RECT  6.420 1.730 6.540 1.900 ;
        RECT  6.405 0.780 6.440 1.195 ;
        RECT  5.670 1.730 6.420 1.850 ;
        RECT  6.230 0.780 6.405 1.555 ;
        RECT  5.760 0.780 6.230 0.900 ;
        RECT  5.910 1.435 6.230 1.555 ;
        RECT  5.790 1.350 5.910 1.610 ;
        RECT  5.550 1.500 5.670 1.850 ;
        RECT  4.920 0.780 5.640 0.900 ;
        RECT  4.920 1.500 5.550 1.620 ;
        RECT  5.310 1.740 5.430 2.140 ;
        RECT  4.005 1.740 5.310 1.860 ;
        RECT  4.800 0.780 4.920 1.620 ;
        RECT  4.620 0.780 4.800 0.900 ;
        RECT  4.620 1.500 4.800 1.620 ;
        RECT  3.960 0.780 4.120 0.900 ;
        RECT  3.960 1.470 4.120 1.590 ;
        RECT  3.885 1.740 4.005 2.100 ;
        RECT  3.870 0.380 3.990 0.655 ;
        RECT  3.840 0.780 3.960 1.590 ;
        RECT  2.440 1.980 3.885 2.100 ;
        RECT  3.480 0.380 3.870 0.500 ;
        RECT  3.600 0.620 3.720 1.860 ;
        RECT  3.010 1.740 3.600 1.860 ;
        RECT  3.360 0.380 3.480 1.620 ;
        RECT  3.155 0.380 3.360 0.810 ;
        RECT  2.890 1.590 3.010 1.860 ;
        RECT  2.340 1.590 2.890 1.710 ;
        RECT  2.580 1.350 2.770 1.470 ;
        RECT  2.460 0.380 2.580 1.470 ;
        RECT  1.610 0.380 2.460 0.500 ;
        RECT  2.320 1.830 2.440 2.100 ;
        RECT  2.220 0.630 2.340 1.710 ;
        RECT  2.020 1.830 2.320 1.950 ;
        RECT  1.820 0.630 2.220 0.750 ;
        RECT  2.130 1.590 2.220 1.710 ;
        RECT  1.800 2.070 2.200 2.190 ;
        RECT  1.980 1.120 2.100 1.470 ;
        RECT  1.900 1.760 2.020 1.950 ;
        RECT  1.385 1.350 1.980 1.470 ;
        RECT  0.600 1.760 1.900 1.880 ;
        RECT  1.680 2.020 1.800 2.190 ;
        RECT  1.210 2.020 1.680 2.140 ;
        RECT  1.490 0.380 1.610 1.210 ;
        RECT  1.080 1.090 1.490 1.210 ;
        RECT  1.265 1.350 1.385 1.540 ;
        RECT  1.020 1.420 1.265 1.540 ;
        RECT  0.950 2.020 1.210 2.150 ;
        RECT  0.960 1.015 1.080 1.275 ;
        RECT  0.840 1.420 1.020 1.620 ;
        RECT  0.840 0.390 0.975 0.895 ;
        RECT  0.805 0.390 0.840 1.620 ;
        RECT  0.760 0.775 0.805 1.620 ;
        RECT  0.720 0.775 0.760 1.540 ;
        RECT  0.480 0.790 0.600 1.880 ;
        RECT  0.255 0.790 0.480 0.910 ;
        RECT  0.255 1.760 0.480 1.880 ;
        RECT  0.085 0.395 0.255 0.910 ;
        RECT  0.085 1.595 0.255 2.025 ;
    END
END AFCSHCONX4AD
MACRO AFCSIHCONX2AD
    CLASS CORE ;
    FOREIGN AFCSIHCONX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.030 0.750 6.090 1.635 ;
        RECT  5.950 0.370 6.030 2.060 ;
        RECT  5.890 0.370 5.950 0.890 ;
        RECT  5.890 1.495 5.950 2.060 ;
        END
        AntennaDiffArea 0.373 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 1.020 5.530 1.655 ;
        END
        AntennaGateArea 0.1817 ;
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.825 1.690 0.875 2.120 ;
        RECT  0.705 1.365 0.825 2.120 ;
        RECT  0.210 1.365 0.705 1.485 ;
        RECT  0.480 0.465 0.600 0.775 ;
        RECT  0.210 0.655 0.480 0.775 ;
        RECT  0.070 0.655 0.210 1.485 ;
        END
        AntennaDiffArea 0.338 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.405 1.485 1.610 2.085 ;
        RECT  1.080 1.485 1.405 1.605 ;
        RECT  1.080 0.750 1.300 0.870 ;
        RECT  0.960 0.750 1.080 1.605 ;
        END
        AntennaDiffArea 0.31 ;
    END CO0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 0.955 1.765 1.125 ;
        RECT  1.490 0.510 1.610 1.125 ;
        RECT  0.840 0.510 1.490 0.630 ;
        RECT  0.720 0.510 0.840 1.065 ;
        RECT  0.335 0.895 0.720 1.065 ;
        END
        AntennaGateArea 0.4408 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 0.940 2.070 1.365 ;
        RECT  1.890 1.245 1.950 1.365 ;
        RECT  1.750 1.245 1.890 1.655 ;
        RECT  1.370 1.245 1.750 1.365 ;
        RECT  1.200 1.030 1.370 1.365 ;
        END
        AntennaGateArea 0.4095 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.685 -0.210 6.160 0.210 ;
        RECT  5.515 -0.210 5.685 0.845 ;
        RECT  4.050 -0.210 5.515 0.210 ;
        RECT  3.880 -0.210 4.050 0.465 ;
        RECT  3.320 -0.210 3.880 0.210 ;
        RECT  3.200 -0.210 3.320 0.880 ;
        RECT  1.955 -0.210 3.200 0.210 ;
        RECT  1.785 -0.210 1.955 0.815 ;
        RECT  1.050 -0.210 1.785 0.210 ;
        RECT  0.790 -0.210 1.050 0.390 ;
        RECT  0.265 -0.210 0.790 0.210 ;
        RECT  0.095 -0.210 0.265 0.535 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.730 2.310 6.160 2.730 ;
        RECT  5.470 2.020 5.730 2.730 ;
        RECT  3.970 2.310 5.470 2.730 ;
        RECT  3.710 1.935 3.970 2.730 ;
        RECT  3.420 2.310 3.710 2.730 ;
        RECT  3.160 1.935 3.420 2.730 ;
        RECT  1.935 2.310 3.160 2.730 ;
        RECT  1.765 1.775 1.935 2.730 ;
        RECT  1.215 2.310 1.765 2.730 ;
        RECT  1.045 1.725 1.215 2.730 ;
        RECT  0.265 2.310 1.045 2.730 ;
        RECT  0.095 1.605 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.770 1.015 5.810 1.275 ;
        RECT  5.650 1.015 5.770 1.900 ;
        RECT  5.265 1.780 5.650 1.900 ;
        RECT  5.150 0.610 5.270 1.640 ;
        RECT  5.145 1.780 5.265 2.125 ;
        RECT  5.050 0.980 5.150 1.240 ;
        RECT  4.595 2.005 5.145 2.125 ;
        RECT  4.920 0.330 5.070 0.450 ;
        RECT  4.920 1.410 4.955 1.840 ;
        RECT  4.810 0.330 4.920 1.840 ;
        RECT  4.785 0.380 4.810 1.840 ;
        RECT  4.290 0.380 4.785 0.500 ;
        RECT  4.595 0.635 4.660 0.805 ;
        RECT  4.410 0.635 4.595 2.125 ;
        RECT  4.170 0.380 4.290 1.090 ;
        RECT  4.115 0.970 4.170 1.090 ;
        RECT  3.940 0.970 4.115 1.795 ;
        RECT  2.675 1.675 3.940 1.795 ;
        RECT  3.535 0.665 3.705 1.505 ;
        RECT  2.840 1.385 3.535 1.505 ;
        RECT  3.080 1.000 3.170 1.260 ;
        RECT  2.960 0.380 3.080 1.260 ;
        RECT  2.315 0.380 2.960 0.500 ;
        RECT  2.720 0.965 2.840 1.505 ;
        RECT  2.600 0.620 2.675 0.790 ;
        RECT  2.600 1.675 2.675 1.860 ;
        RECT  2.480 0.620 2.600 1.860 ;
        RECT  2.190 0.365 2.315 1.920 ;
        RECT  2.145 0.365 2.190 0.795 ;
        RECT  2.145 1.490 2.190 1.920 ;
    END
END AFCSIHCONX2AD
MACRO AFCSIHCONX4AD
    CLASS CORE ;
    FOREIGN AFCSIHCONX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.465 1.005 7.490 1.515 ;
        RECT  7.345 0.370 7.465 2.030 ;
        RECT  7.300 0.370 7.345 0.890 ;
        RECT  7.300 1.510 7.345 2.030 ;
        END
        AntennaDiffArea 0.373 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.710 1.030 6.930 1.375 ;
        END
        AntennaGateArea 0.1825 ;
    END CS
    PIN CO1N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.315 1.495 1.485 1.670 ;
        RECT  1.215 0.515 1.385 0.750 ;
        RECT  0.240 1.495 1.315 1.625 ;
        RECT  0.665 0.620 1.215 0.750 ;
        RECT  0.495 0.515 0.665 0.750 ;
        RECT  0.210 0.620 0.495 0.750 ;
        RECT  0.210 1.495 0.240 2.085 ;
        RECT  0.070 0.620 0.210 2.085 ;
        END
        AntennaDiffArea 0.666 ;
    END CO1N
    PIN CO0N
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.675 1.470 2.845 2.005 ;
        RECT  2.255 1.470 2.675 1.610 ;
        RECT  2.255 0.675 2.465 0.795 ;
        RECT  2.125 0.675 2.255 1.610 ;
        RECT  2.115 0.675 2.125 1.975 ;
        RECT  1.955 1.470 2.115 1.975 ;
        END
        AntennaDiffArea 0.559 ;
    END CO0N
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.770 0.990 2.955 1.110 ;
        RECT  2.650 0.420 2.770 1.110 ;
        RECT  1.990 0.420 2.650 0.540 ;
        RECT  1.870 0.420 1.990 1.235 ;
        RECT  1.820 0.975 1.870 1.235 ;
        RECT  1.700 0.975 1.820 1.330 ;
        RECT  0.970 1.190 1.700 1.330 ;
        RECT  0.710 1.120 0.970 1.330 ;
        END
        AntennaGateArea 0.7298 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.955 3.290 1.655 ;
        RECT  2.530 1.230 3.150 1.350 ;
        RECT  2.380 1.060 2.530 1.350 ;
        END
        AntennaGateArea 0.6962 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.130 -0.210 7.560 0.210 ;
        RECT  6.870 -0.210 7.130 0.690 ;
        RECT  5.305 -0.210 6.870 0.210 ;
        RECT  5.135 -0.210 5.305 0.740 ;
        RECT  4.580 -0.210 5.135 0.210 ;
        RECT  4.440 -0.210 4.580 0.900 ;
        RECT  3.060 -0.210 4.440 0.210 ;
        RECT  2.890 -0.210 3.060 0.725 ;
        RECT  1.750 -0.210 2.890 0.210 ;
        RECT  1.580 -0.210 1.750 0.720 ;
        RECT  1.025 -0.210 1.580 0.210 ;
        RECT  0.855 -0.210 1.025 0.490 ;
        RECT  0.305 -0.210 0.855 0.210 ;
        RECT  0.135 -0.210 0.305 0.490 ;
        RECT  0.000 -0.210 0.135 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.085 2.310 7.560 2.730 ;
        RECT  6.915 1.980 7.085 2.730 ;
        RECT  5.330 2.310 6.915 2.730 ;
        RECT  5.070 2.105 5.330 2.730 ;
        RECT  4.680 2.310 5.070 2.730 ;
        RECT  4.420 2.105 4.680 2.730 ;
        RECT  3.205 2.310 4.420 2.730 ;
        RECT  3.035 1.775 3.205 2.730 ;
        RECT  2.485 2.310 3.035 2.730 ;
        RECT  2.315 1.735 2.485 2.730 ;
        RECT  1.765 2.310 2.315 2.730 ;
        RECT  1.595 1.830 1.765 2.730 ;
        RECT  0.920 2.310 1.595 2.730 ;
        RECT  0.660 1.745 0.920 2.730 ;
        RECT  0.000 2.310 0.660 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  7.170 1.015 7.225 1.275 ;
        RECT  7.050 1.015 7.170 1.855 ;
        RECT  6.745 1.735 7.050 1.855 ;
        RECT  6.530 1.495 6.750 1.615 ;
        RECT  6.575 1.735 6.745 2.140 ;
        RECT  6.560 0.505 6.680 0.910 ;
        RECT  5.925 2.020 6.575 2.140 ;
        RECT  6.530 0.790 6.560 0.910 ;
        RECT  6.410 0.790 6.530 1.615 ;
        RECT  6.105 0.335 6.275 1.900 ;
        RECT  5.545 0.380 6.105 0.500 ;
        RECT  5.925 0.620 5.960 0.740 ;
        RECT  5.745 0.620 5.925 2.140 ;
        RECT  5.700 0.620 5.745 0.740 ;
        RECT  5.425 0.380 5.545 1.250 ;
        RECT  5.195 1.080 5.425 1.250 ;
        RECT  5.070 1.080 5.195 1.975 ;
        RECT  3.810 1.855 5.070 1.975 ;
        RECT  4.830 0.640 4.950 1.655 ;
        RECT  4.820 0.640 4.830 1.480 ;
        RECT  4.050 1.360 4.820 1.480 ;
        RECT  4.320 1.035 4.415 1.215 ;
        RECT  4.200 0.380 4.320 1.215 ;
        RECT  3.540 0.380 4.200 0.500 ;
        RECT  3.930 0.980 4.050 1.480 ;
        RECT  3.810 0.620 3.865 0.790 ;
        RECT  3.690 0.620 3.810 1.975 ;
        RECT  3.420 0.380 3.540 1.940 ;
        RECT  3.275 0.380 3.420 0.810 ;
        RECT  1.335 0.870 1.505 1.045 ;
        RECT  0.330 0.870 1.335 0.990 ;
    END
END AFCSIHCONX4AD
MACRO AFHCINX2AD
    CLASS CORE ;
    FOREIGN AFHCINX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.630 0.670 7.770 1.760 ;
        RECT  7.380 0.670 7.630 0.790 ;
        RECT  7.430 1.500 7.630 1.760 ;
        END
        AntennaDiffArea 0.251 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.385 1.450 5.505 1.880 ;
        RECT  4.785 1.760 5.385 1.880 ;
        RECT  5.020 0.525 5.170 0.955 ;
        RECT  4.900 0.525 5.020 1.330 ;
        RECT  4.785 1.190 4.900 1.330 ;
        RECT  4.665 1.190 4.785 1.880 ;
        END
        AntennaDiffArea 0.518 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.800 1.145 8.890 1.375 ;
        RECT  8.615 0.995 8.800 1.375 ;
        END
        AntennaGateArea 0.3204 ;
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.595 0.950 3.715 1.260 ;
        RECT  3.570 0.950 3.595 1.070 ;
        RECT  3.450 0.750 3.570 1.070 ;
        RECT  3.335 0.750 3.450 0.870 ;
        RECT  3.210 0.350 3.335 0.870 ;
        RECT  3.105 0.350 3.210 0.490 ;
        END
        AntennaGateArea 0.4454 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.055 0.400 1.225 ;
        RECT  0.070 0.880 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.875 -0.210 8.960 0.210 ;
        RECT  8.705 -0.210 8.875 0.845 ;
        RECT  7.910 -0.210 8.705 0.210 ;
        RECT  7.650 -0.210 7.910 0.230 ;
        RECT  7.260 -0.210 7.650 0.210 ;
        RECT  7.000 -0.210 7.260 0.230 ;
        RECT  4.060 -0.210 7.000 0.210 ;
        RECT  3.800 -0.210 4.060 0.390 ;
        RECT  0.875 -0.210 3.800 0.210 ;
        RECT  0.445 -0.210 0.875 0.415 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.875 2.310 8.960 2.730 ;
        RECT  8.705 1.575 8.875 2.730 ;
        RECT  7.740 2.310 8.705 2.730 ;
        RECT  7.220 2.270 7.740 2.730 ;
        RECT  3.920 2.310 7.220 2.730 ;
        RECT  3.660 2.290 3.920 2.730 ;
        RECT  0.660 2.310 3.660 2.730 ;
        RECT  0.400 2.010 0.660 2.730 ;
        RECT  0.000 2.310 0.400 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.960 2.520 ;
        LAYER M1 ;
        RECT  8.370 0.350 8.490 2.090 ;
        RECT  7.290 1.970 8.370 2.090 ;
        RECT  8.100 0.380 8.220 1.745 ;
        RECT  5.505 0.380 8.100 0.500 ;
        RECT  7.380 0.940 7.500 1.250 ;
        RECT  7.150 0.940 7.380 1.060 ;
        RECT  7.170 1.350 7.290 2.090 ;
        RECT  7.100 1.350 7.170 1.470 ;
        RECT  6.950 1.970 7.170 2.090 ;
        RECT  7.030 0.620 7.150 1.060 ;
        RECT  6.980 1.180 7.100 1.470 ;
        RECT  6.420 0.620 7.030 0.740 ;
        RECT  6.845 1.970 6.950 2.140 ;
        RECT  6.855 1.615 6.905 1.785 ;
        RECT  6.855 0.860 6.880 0.980 ;
        RECT  6.735 0.860 6.855 1.785 ;
        RECT  6.185 2.020 6.845 2.140 ;
        RECT  6.620 0.860 6.735 0.980 ;
        RECT  6.495 1.725 6.545 1.895 ;
        RECT  6.420 1.195 6.495 1.895 ;
        RECT  6.375 0.620 6.420 1.895 ;
        RECT  6.300 0.620 6.375 1.315 ;
        RECT  5.745 0.620 6.300 0.740 ;
        RECT  6.135 1.725 6.185 2.140 ;
        RECT  6.015 0.860 6.135 2.140 ;
        RECT  5.875 0.860 6.015 1.030 ;
        RECT  5.745 1.220 5.775 2.050 ;
        RECT  5.655 0.620 5.745 2.050 ;
        RECT  5.625 0.620 5.655 1.340 ;
        RECT  5.385 0.380 5.505 1.220 ;
        RECT  5.195 2.020 5.455 2.180 ;
        RECT  5.265 1.090 5.385 1.220 ;
        RECT  5.145 1.090 5.265 1.640 ;
        RECT  2.610 2.020 5.195 2.140 ;
        RECT  4.955 1.520 5.145 1.640 ;
        RECT  4.660 0.475 4.780 0.735 ;
        RECT  4.375 0.615 4.660 0.735 ;
        RECT  4.425 0.880 4.545 1.900 ;
        RECT  2.850 1.780 4.425 1.900 ;
        RECT  4.300 0.540 4.375 0.735 ;
        RECT  4.180 0.540 4.300 1.660 ;
        RECT  4.160 1.400 4.180 1.660 ;
        RECT  4.015 1.005 4.060 1.265 ;
        RECT  3.895 0.510 4.015 1.560 ;
        RECT  3.590 0.510 3.895 0.630 ;
        RECT  3.575 1.440 3.895 1.560 ;
        RECT  3.470 0.370 3.590 0.630 ;
        RECT  3.475 1.440 3.575 1.610 ;
        RECT  3.405 1.205 3.475 1.610 ;
        RECT  3.355 1.205 3.405 1.560 ;
        RECT  3.330 1.205 3.355 1.325 ;
        RECT  3.210 0.990 3.330 1.325 ;
        RECT  3.090 1.485 3.235 1.655 ;
        RECT  2.970 0.650 3.090 1.655 ;
        RECT  2.895 0.650 2.970 0.770 ;
        RECT  2.725 0.380 2.895 0.770 ;
        RECT  2.730 0.890 2.850 1.900 ;
        RECT  2.510 0.890 2.730 1.010 ;
        RECT  1.210 0.380 2.725 0.500 ;
        RECT  2.490 1.130 2.610 2.140 ;
        RECT  2.390 0.625 2.510 1.010 ;
        RECT  2.270 1.130 2.490 1.250 ;
        RECT  2.100 2.020 2.490 2.140 ;
        RECT  2.250 1.370 2.370 1.825 ;
        RECT  2.150 0.620 2.270 1.250 ;
        RECT  1.860 1.370 2.250 1.490 ;
        RECT  1.500 0.620 2.150 0.740 ;
        RECT  1.970 1.715 2.100 2.140 ;
        RECT  1.860 0.870 2.000 0.990 ;
        RECT  1.840 1.715 1.970 1.835 ;
        RECT  1.740 0.870 1.860 1.490 ;
        RECT  1.670 1.370 1.740 1.490 ;
        RECT  1.550 1.370 1.670 2.140 ;
        RECT  0.910 2.020 1.550 2.140 ;
        RECT  1.380 0.620 1.500 1.195 ;
        RECT  1.335 1.075 1.380 1.195 ;
        RECT  1.215 1.075 1.335 1.900 ;
        RECT  1.165 1.730 1.215 1.900 ;
        RECT  1.090 0.380 1.210 0.905 ;
        RECT  1.070 0.785 1.090 0.905 ;
        RECT  0.950 0.785 1.070 1.650 ;
        RECT  0.760 1.530 0.950 1.650 ;
        RECT  0.790 1.770 0.910 2.140 ;
        RECT  0.645 0.970 0.830 1.230 ;
        RECT  0.640 1.770 0.790 1.890 ;
        RECT  0.640 0.640 0.645 1.230 ;
        RECT  0.520 0.640 0.640 1.890 ;
        RECT  0.255 0.640 0.520 0.760 ;
        RECT  0.255 1.770 0.520 1.890 ;
        RECT  0.085 0.330 0.255 0.760 ;
        RECT  0.085 1.600 0.255 2.030 ;
    END
END AFHCINX2AD
MACRO AFHCINX4AD
    CLASS CORE ;
    FOREIGN AFHCINX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.590 0.670 9.730 1.715 ;
        RECT  9.400 0.670 9.590 0.790 ;
        RECT  9.425 1.545 9.590 1.715 ;
        END
        AntennaDiffArea 0.254 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.210 0.665 7.295 0.835 ;
        RECT  7.155 0.665 7.210 1.400 ;
        RECT  7.070 0.665 7.155 1.900 ;
        RECT  7.030 1.235 7.070 1.900 ;
        RECT  5.625 1.780 7.030 1.900 ;
        RECT  6.405 0.525 6.575 0.955 ;
        RECT  6.400 0.525 6.405 0.910 ;
        RECT  5.625 0.790 6.400 0.910 ;
        RECT  5.505 0.790 5.625 1.900 ;
        RECT  4.715 1.780 5.505 1.900 ;
        END
        AntennaDiffArea 1.037 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.570 1.065 10.865 1.235 ;
        RECT  10.430 1.065 10.570 1.375 ;
        END
        AntennaGateArea 0.648 ;
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.990 1.000 4.155 1.375 ;
        END
        AntennaGateArea 0.4787 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.055 0.375 1.225 ;
        RECT  0.070 0.880 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.395 -0.210 11.480 0.210 ;
        RECT  11.225 -0.210 11.395 0.675 ;
        RECT  10.675 -0.210 11.225 0.210 ;
        RECT  10.505 -0.210 10.675 0.675 ;
        RECT  9.930 -0.210 10.505 0.210 ;
        RECT  9.670 -0.210 9.930 0.230 ;
        RECT  9.230 -0.210 9.670 0.210 ;
        RECT  8.970 -0.210 9.230 0.230 ;
        RECT  4.485 -0.210 8.970 0.210 ;
        RECT  4.225 -0.210 4.485 0.390 ;
        RECT  0.875 -0.210 4.225 0.210 ;
        RECT  0.445 -0.210 0.875 0.415 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.395 2.310 11.480 2.730 ;
        RECT  11.225 1.845 11.395 2.730 ;
        RECT  10.675 2.310 11.225 2.730 ;
        RECT  10.505 2.085 10.675 2.730 ;
        RECT  9.915 2.310 10.505 2.730 ;
        RECT  9.135 2.260 9.915 2.730 ;
        RECT  4.300 2.310 9.135 2.730 ;
        RECT  4.130 2.105 4.300 2.730 ;
        RECT  0.660 2.310 4.130 2.730 ;
        RECT  0.400 2.010 0.660 2.730 ;
        RECT  0.000 2.310 0.400 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.480 2.520 ;
        LAYER M1 ;
        RECT  11.010 0.810 11.110 1.590 ;
        RECT  10.990 0.410 11.010 1.955 ;
        RECT  10.890 0.410 10.990 0.930 ;
        RECT  10.890 1.435 10.990 1.955 ;
        RECT  9.130 1.835 10.890 1.955 ;
        RECT  10.170 0.380 10.290 1.590 ;
        RECT  6.910 0.380 10.170 0.500 ;
        RECT  9.300 0.940 9.420 1.320 ;
        RECT  9.120 0.940 9.300 1.060 ;
        RECT  9.070 1.350 9.130 2.090 ;
        RECT  9.000 0.620 9.120 1.060 ;
        RECT  9.010 1.180 9.070 2.090 ;
        RECT  8.950 1.180 9.010 1.470 ;
        RECT  8.910 1.970 9.010 2.090 ;
        RECT  8.420 0.620 9.000 0.740 ;
        RECT  8.805 1.970 8.910 2.140 ;
        RECT  8.825 1.615 8.875 1.785 ;
        RECT  8.825 0.860 8.850 0.980 ;
        RECT  8.705 0.860 8.825 1.785 ;
        RECT  8.155 2.020 8.805 2.140 ;
        RECT  8.590 0.860 8.705 0.980 ;
        RECT  8.465 1.725 8.515 1.895 ;
        RECT  8.420 1.195 8.465 1.895 ;
        RECT  8.345 0.620 8.420 1.895 ;
        RECT  8.300 0.620 8.345 1.315 ;
        RECT  7.635 0.620 8.300 0.740 ;
        RECT  8.105 1.725 8.155 2.140 ;
        RECT  7.985 0.860 8.105 2.140 ;
        RECT  7.800 0.860 7.985 0.980 ;
        RECT  7.410 2.020 7.985 2.140 ;
        RECT  7.650 1.220 7.770 1.750 ;
        RECT  7.635 1.220 7.650 1.340 ;
        RECT  7.515 0.620 7.635 1.340 ;
        RECT  7.465 0.620 7.515 0.790 ;
        RECT  7.290 1.680 7.410 2.140 ;
        RECT  6.790 0.380 6.910 1.640 ;
        RECT  6.600 2.020 6.860 2.180 ;
        RECT  6.105 1.230 6.790 1.360 ;
        RECT  6.515 1.520 6.790 1.640 ;
        RECT  6.395 2.020 6.600 2.140 ;
        RECT  6.135 2.020 6.395 2.180 ;
        RECT  5.385 0.550 6.260 0.670 ;
        RECT  5.935 2.020 6.135 2.140 ;
        RECT  5.985 1.230 6.105 1.640 ;
        RECT  5.795 1.520 5.985 1.640 ;
        RECT  5.675 2.020 5.935 2.180 ;
        RECT  4.550 2.020 5.675 2.140 ;
        RECT  5.265 0.380 5.385 1.640 ;
        RECT  4.605 0.380 5.265 0.500 ;
        RECT  4.635 1.520 5.265 1.640 ;
        RECT  4.995 0.620 5.115 1.320 ;
        RECT  4.485 0.620 4.995 0.740 ;
        RECT  4.515 1.330 4.635 1.640 ;
        RECT  4.395 1.075 4.585 1.195 ;
        RECT  4.430 1.805 4.550 2.140 ;
        RECT  4.365 0.510 4.485 0.740 ;
        RECT  4.000 1.805 4.430 1.925 ;
        RECT  4.275 1.075 4.395 1.620 ;
        RECT  3.565 0.510 4.365 0.630 ;
        RECT  3.805 1.500 4.275 1.620 ;
        RECT  3.805 0.760 4.105 0.880 ;
        RECT  3.880 1.805 4.000 2.070 ;
        RECT  2.675 1.950 3.880 2.070 ;
        RECT  3.685 0.760 3.805 1.620 ;
        RECT  3.445 0.510 3.565 1.830 ;
        RECT  2.990 1.710 3.445 1.830 ;
        RECT  3.205 0.380 3.325 1.590 ;
        RECT  3.180 0.380 3.205 0.740 ;
        RECT  1.210 0.380 3.180 0.500 ;
        RECT  2.965 1.400 2.990 1.830 ;
        RECT  2.845 0.675 2.965 1.830 ;
        RECT  2.535 0.675 2.845 0.845 ;
        RECT  2.820 1.400 2.845 1.830 ;
        RECT  2.555 1.715 2.675 2.070 ;
        RECT  2.410 1.715 2.555 1.835 ;
        RECT  2.265 1.970 2.435 2.140 ;
        RECT  2.290 0.620 2.410 1.835 ;
        RECT  1.500 0.620 2.290 0.740 ;
        RECT  2.055 1.715 2.290 1.835 ;
        RECT  1.670 2.020 2.265 2.140 ;
        RECT  1.885 0.860 2.115 0.980 ;
        RECT  1.885 1.715 2.055 1.885 ;
        RECT  1.765 0.860 1.885 1.585 ;
        RECT  1.670 1.465 1.765 1.585 ;
        RECT  1.550 1.465 1.670 2.140 ;
        RECT  0.910 2.020 1.550 2.140 ;
        RECT  1.380 0.620 1.500 1.325 ;
        RECT  1.335 1.205 1.380 1.325 ;
        RECT  1.215 1.205 1.335 1.900 ;
        RECT  1.165 1.730 1.215 1.900 ;
        RECT  1.090 0.380 1.210 1.010 ;
        RECT  1.020 0.890 1.090 1.010 ;
        RECT  0.900 0.890 1.020 1.650 ;
        RECT  0.790 1.770 0.910 2.140 ;
        RECT  0.760 1.530 0.900 1.650 ;
        RECT  0.640 1.770 0.790 1.890 ;
        RECT  0.645 0.970 0.715 1.230 ;
        RECT  0.640 0.640 0.645 1.230 ;
        RECT  0.520 0.640 0.640 1.890 ;
        RECT  0.255 0.640 0.520 0.760 ;
        RECT  0.255 1.770 0.520 1.890 ;
        RECT  0.085 0.330 0.255 0.760 ;
        RECT  0.085 1.600 0.255 2.030 ;
    END
END AFHCINX4AD
MACRO AFHCONX2AD
    CLASS CORE ;
    FOREIGN AFHCONX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.630 0.670 7.770 1.760 ;
        RECT  7.380 0.670 7.630 0.790 ;
        RECT  7.430 1.500 7.630 1.760 ;
        END
        AntennaDiffArea 0.251 ;
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.410 1.465 5.530 1.880 ;
        RECT  4.800 1.760 5.410 1.880 ;
        RECT  5.050 0.525 5.195 0.955 ;
        RECT  4.930 0.525 5.050 1.330 ;
        RECT  4.800 1.190 4.930 1.330 ;
        RECT  4.680 1.190 4.800 1.880 ;
        END
        AntennaDiffArea 0.504 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.800 1.145 8.890 1.375 ;
        RECT  8.615 0.995 8.800 1.375 ;
        END
        AntennaGateArea 0.3184 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.655 1.000 3.775 1.260 ;
        RECT  3.570 1.000 3.655 1.120 ;
        RECT  3.450 0.800 3.570 1.120 ;
        RECT  3.335 0.800 3.450 0.920 ;
        RECT  3.210 0.350 3.335 0.920 ;
        RECT  3.105 0.350 3.210 0.490 ;
        END
        AntennaGateArea 0.4989 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.055 0.400 1.225 ;
        RECT  0.070 0.880 0.210 1.375 ;
        END
        AntennaGateArea 0.16 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.875 -0.210 8.960 0.210 ;
        RECT  8.705 -0.210 8.875 0.845 ;
        RECT  7.910 -0.210 8.705 0.210 ;
        RECT  7.650 -0.210 7.910 0.230 ;
        RECT  7.260 -0.210 7.650 0.210 ;
        RECT  7.000 -0.210 7.260 0.230 ;
        RECT  4.060 -0.210 7.000 0.210 ;
        RECT  3.800 -0.210 4.060 0.390 ;
        RECT  0.875 -0.210 3.800 0.210 ;
        RECT  0.445 -0.210 0.875 0.435 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.875 2.310 8.960 2.730 ;
        RECT  8.705 1.575 8.875 2.730 ;
        RECT  7.740 2.310 8.705 2.730 ;
        RECT  7.220 2.270 7.740 2.730 ;
        RECT  3.920 2.310 7.220 2.730 ;
        RECT  3.660 2.290 3.920 2.730 ;
        RECT  0.660 2.310 3.660 2.730 ;
        RECT  0.400 2.010 0.660 2.730 ;
        RECT  0.000 2.310 0.400 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.960 2.520 ;
        LAYER M1 ;
        RECT  8.370 0.350 8.490 2.090 ;
        RECT  7.290 1.970 8.370 2.090 ;
        RECT  8.100 0.380 8.220 1.745 ;
        RECT  5.530 0.380 8.100 0.500 ;
        RECT  7.380 0.940 7.500 1.250 ;
        RECT  7.150 0.940 7.380 1.060 ;
        RECT  7.170 1.350 7.290 2.090 ;
        RECT  7.100 1.350 7.170 1.470 ;
        RECT  6.950 1.970 7.170 2.090 ;
        RECT  7.030 0.620 7.150 1.060 ;
        RECT  6.980 1.180 7.100 1.470 ;
        RECT  6.420 0.620 7.030 0.740 ;
        RECT  6.845 1.970 6.950 2.140 ;
        RECT  6.855 1.615 6.905 1.785 ;
        RECT  6.855 0.860 6.880 0.980 ;
        RECT  6.735 0.860 6.855 1.785 ;
        RECT  6.185 2.020 6.845 2.140 ;
        RECT  6.620 0.860 6.735 0.980 ;
        RECT  6.495 1.780 6.590 1.900 ;
        RECT  6.420 1.195 6.495 1.900 ;
        RECT  6.375 0.620 6.420 1.900 ;
        RECT  6.300 0.620 6.375 1.315 ;
        RECT  6.330 1.780 6.375 1.900 ;
        RECT  5.770 0.620 6.300 0.740 ;
        RECT  6.135 1.830 6.185 2.140 ;
        RECT  6.015 0.860 6.135 2.140 ;
        RECT  5.895 0.860 6.015 1.030 ;
        RECT  5.770 1.220 5.800 2.145 ;
        RECT  5.680 0.620 5.770 2.145 ;
        RECT  5.650 0.620 5.680 1.340 ;
        RECT  5.410 0.380 5.530 1.220 ;
        RECT  5.290 1.090 5.410 1.220 ;
        RECT  4.380 2.020 5.380 2.140 ;
        RECT  5.170 1.090 5.290 1.640 ;
        RECT  4.980 1.520 5.170 1.640 ;
        RECT  4.690 0.470 4.810 0.730 ;
        RECT  4.375 0.610 4.690 0.730 ;
        RECT  4.440 0.850 4.560 1.870 ;
        RECT  2.850 1.750 4.440 1.870 ;
        RECT  4.260 1.990 4.380 2.140 ;
        RECT  4.280 0.540 4.375 0.730 ;
        RECT  4.160 0.540 4.280 1.620 ;
        RECT  2.610 1.990 4.260 2.110 ;
        RECT  3.895 0.560 4.015 1.560 ;
        RECT  3.590 0.560 3.895 0.680 ;
        RECT  3.575 1.440 3.895 1.560 ;
        RECT  3.470 0.420 3.590 0.680 ;
        RECT  3.525 1.440 3.575 1.610 ;
        RECT  3.405 1.255 3.525 1.610 ;
        RECT  3.330 1.255 3.405 1.375 ;
        RECT  3.210 1.045 3.330 1.375 ;
        RECT  3.090 1.510 3.280 1.630 ;
        RECT  2.970 0.650 3.090 1.630 ;
        RECT  2.895 0.650 2.970 0.770 ;
        RECT  2.725 0.380 2.895 0.770 ;
        RECT  2.730 0.890 2.850 1.870 ;
        RECT  2.510 0.890 2.730 1.010 ;
        RECT  1.210 0.380 2.725 0.500 ;
        RECT  2.490 1.130 2.610 2.110 ;
        RECT  2.390 0.625 2.510 1.010 ;
        RECT  2.270 1.130 2.490 1.250 ;
        RECT  2.100 1.990 2.490 2.110 ;
        RECT  2.250 1.370 2.370 1.825 ;
        RECT  2.150 0.620 2.270 1.250 ;
        RECT  1.860 1.370 2.250 1.490 ;
        RECT  1.500 0.620 2.150 0.740 ;
        RECT  1.970 1.715 2.100 2.110 ;
        RECT  1.860 0.870 2.000 0.990 ;
        RECT  1.840 1.715 1.970 1.835 ;
        RECT  1.740 0.870 1.860 1.490 ;
        RECT  1.670 1.370 1.740 1.490 ;
        RECT  1.550 1.370 1.670 2.140 ;
        RECT  0.910 2.020 1.550 2.140 ;
        RECT  1.380 0.620 1.500 1.195 ;
        RECT  1.335 1.075 1.380 1.195 ;
        RECT  1.215 1.075 1.335 1.900 ;
        RECT  1.165 1.730 1.215 1.900 ;
        RECT  1.090 0.380 1.210 0.905 ;
        RECT  1.070 0.785 1.090 0.905 ;
        RECT  0.950 0.785 1.070 1.650 ;
        RECT  0.760 1.530 0.950 1.650 ;
        RECT  0.790 1.770 0.910 2.140 ;
        RECT  0.645 0.970 0.830 1.230 ;
        RECT  0.640 1.770 0.790 1.890 ;
        RECT  0.640 0.640 0.645 1.230 ;
        RECT  0.520 0.640 0.640 1.890 ;
        RECT  0.255 0.640 0.520 0.760 ;
        RECT  0.255 1.770 0.520 1.890 ;
        RECT  0.085 0.330 0.255 0.760 ;
        RECT  0.085 1.600 0.255 2.030 ;
    END
END AFHCONX2AD
MACRO AFHCONX4AD
    CLASS CORE ;
    FOREIGN AFHCONX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.190 0.670 8.330 1.760 ;
        RECT  7.850 0.670 8.190 0.790 ;
        RECT  7.850 1.500 8.190 1.760 ;
        END
        AntennaDiffArea 0.251 ;
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.810 0.620 5.860 1.055 ;
        RECT  5.740 0.620 5.810 1.515 ;
        RECT  5.670 0.935 5.740 1.515 ;
        RECT  5.520 1.395 5.670 1.515 ;
        RECT  5.400 1.395 5.520 1.880 ;
        RECT  4.790 1.760 5.400 1.880 ;
        RECT  5.040 0.655 5.165 0.825 ;
        RECT  4.920 0.655 5.040 1.330 ;
        RECT  4.790 1.190 4.920 1.330 ;
        RECT  4.670 1.190 4.790 1.880 ;
        END
        AntennaDiffArea 0.696 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.985 0.995 9.190 1.375 ;
        RECT  8.810 0.995 8.985 1.255 ;
        END
        AntennaGateArea 0.482 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.655 1.000 3.775 1.260 ;
        RECT  3.570 1.000 3.655 1.120 ;
        RECT  3.450 0.800 3.570 1.120 ;
        RECT  3.335 0.800 3.450 0.920 ;
        RECT  3.210 0.350 3.335 0.920 ;
        RECT  3.105 0.350 3.210 0.490 ;
        END
        AntennaGateArea 0.4989 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.055 0.400 1.225 ;
        RECT  0.070 0.880 0.210 1.375 ;
        END
        AntennaGateArea 0.16 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.075 -0.210 9.520 0.210 ;
        RECT  8.905 -0.210 9.075 0.720 ;
        RECT  8.380 -0.210 8.905 0.210 ;
        RECT  8.120 -0.210 8.380 0.230 ;
        RECT  7.730 -0.210 8.120 0.210 ;
        RECT  7.470 -0.210 7.730 0.230 ;
        RECT  4.060 -0.210 7.470 0.210 ;
        RECT  3.800 -0.210 4.060 0.390 ;
        RECT  0.875 -0.210 3.800 0.210 ;
        RECT  0.445 -0.210 0.875 0.435 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.120 2.310 9.520 2.730 ;
        RECT  8.860 2.130 9.120 2.730 ;
        RECT  8.160 2.310 8.860 2.730 ;
        RECT  7.640 2.270 8.160 2.730 ;
        RECT  3.920 2.310 7.640 2.730 ;
        RECT  3.660 2.290 3.920 2.730 ;
        RECT  0.660 2.310 3.660 2.730 ;
        RECT  0.400 2.010 0.660 2.730 ;
        RECT  0.000 2.310 0.400 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.520 2.520 ;
        LAYER M1 ;
        RECT  9.315 0.435 9.435 2.000 ;
        RECT  9.265 0.435 9.315 0.865 ;
        RECT  9.265 1.570 9.315 2.000 ;
        RECT  7.570 1.880 9.265 2.000 ;
        RECT  8.570 0.380 8.690 1.745 ;
        RECT  6.100 0.380 8.570 0.500 ;
        RECT  7.800 0.940 7.920 1.275 ;
        RECT  7.730 0.940 7.800 1.060 ;
        RECT  7.610 0.620 7.730 1.060 ;
        RECT  7.010 0.620 7.610 0.740 ;
        RECT  7.520 1.270 7.570 2.090 ;
        RECT  7.450 1.180 7.520 2.090 ;
        RECT  7.400 1.180 7.450 1.440 ;
        RECT  7.370 1.970 7.450 2.090 ;
        RECT  7.275 0.860 7.440 0.980 ;
        RECT  7.265 1.970 7.370 2.140 ;
        RECT  7.275 1.575 7.325 1.745 ;
        RECT  7.155 0.860 7.275 1.745 ;
        RECT  6.580 2.020 7.265 2.140 ;
        RECT  6.890 0.620 7.010 1.900 ;
        RECT  6.390 0.620 6.890 0.740 ;
        RECT  6.750 1.780 6.890 1.900 ;
        RECT  6.580 0.860 6.630 1.660 ;
        RECT  6.510 0.860 6.580 2.140 ;
        RECT  6.460 1.540 6.510 2.140 ;
        RECT  6.340 0.620 6.390 1.365 ;
        RECT  6.270 0.620 6.340 2.075 ;
        RECT  6.220 1.245 6.270 2.075 ;
        RECT  6.030 1.955 6.220 2.075 ;
        RECT  5.980 0.380 6.100 1.755 ;
        RECT  5.500 0.380 5.980 0.500 ;
        RECT  5.880 1.635 5.980 1.755 ;
        RECT  5.760 1.635 5.880 1.895 ;
        RECT  5.540 2.020 5.800 2.160 ;
        RECT  2.610 2.020 5.540 2.140 ;
        RECT  5.380 0.380 5.500 1.220 ;
        RECT  5.280 1.090 5.380 1.220 ;
        RECT  5.160 1.090 5.280 1.640 ;
        RECT  4.970 1.520 5.160 1.640 ;
        RECT  4.660 0.470 4.780 0.730 ;
        RECT  4.375 0.610 4.660 0.730 ;
        RECT  4.430 0.850 4.550 1.900 ;
        RECT  2.850 1.780 4.430 1.900 ;
        RECT  4.280 0.540 4.375 0.730 ;
        RECT  4.160 0.540 4.280 1.660 ;
        RECT  3.895 0.560 4.015 1.560 ;
        RECT  3.590 0.560 3.895 0.680 ;
        RECT  3.575 1.440 3.895 1.560 ;
        RECT  3.470 0.420 3.590 0.680 ;
        RECT  3.525 1.440 3.575 1.610 ;
        RECT  3.405 1.255 3.525 1.610 ;
        RECT  3.330 1.255 3.405 1.375 ;
        RECT  3.210 1.045 3.330 1.375 ;
        RECT  3.090 1.510 3.280 1.630 ;
        RECT  2.970 0.650 3.090 1.630 ;
        RECT  2.895 0.650 2.970 0.770 ;
        RECT  2.725 0.380 2.895 0.770 ;
        RECT  2.730 0.890 2.850 1.900 ;
        RECT  2.510 0.890 2.730 1.010 ;
        RECT  1.210 0.380 2.725 0.500 ;
        RECT  2.490 1.130 2.610 2.140 ;
        RECT  2.390 0.625 2.510 1.010 ;
        RECT  2.270 1.130 2.490 1.250 ;
        RECT  2.100 2.020 2.490 2.140 ;
        RECT  2.250 1.370 2.370 1.825 ;
        RECT  2.150 0.620 2.270 1.250 ;
        RECT  1.860 1.370 2.250 1.490 ;
        RECT  1.500 0.620 2.150 0.740 ;
        RECT  1.970 1.715 2.100 2.140 ;
        RECT  1.860 0.870 2.000 0.990 ;
        RECT  1.840 1.715 1.970 1.835 ;
        RECT  1.740 0.870 1.860 1.490 ;
        RECT  1.670 1.370 1.740 1.490 ;
        RECT  1.550 1.370 1.670 2.140 ;
        RECT  0.910 2.020 1.550 2.140 ;
        RECT  1.380 0.620 1.500 1.195 ;
        RECT  1.335 1.075 1.380 1.195 ;
        RECT  1.215 1.075 1.335 1.900 ;
        RECT  1.165 1.730 1.215 1.900 ;
        RECT  1.090 0.380 1.210 0.905 ;
        RECT  1.070 0.785 1.090 0.905 ;
        RECT  0.950 0.785 1.070 1.650 ;
        RECT  0.760 1.530 0.950 1.650 ;
        RECT  0.790 1.770 0.910 2.140 ;
        RECT  0.645 0.970 0.830 1.230 ;
        RECT  0.640 1.770 0.790 1.890 ;
        RECT  0.640 0.640 0.645 1.230 ;
        RECT  0.520 0.640 0.640 1.890 ;
        RECT  0.255 0.640 0.520 0.760 ;
        RECT  0.255 1.770 0.520 1.890 ;
        RECT  0.085 0.330 0.255 0.760 ;
        RECT  0.085 1.600 0.255 2.030 ;
    END
END AFHCONX4AD
MACRO AHCSHCINX2AD
    CLASS CORE ;
    FOREIGN AHCSHCINX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.090 0.400 5.250 1.965 ;
        END
        AntennaDiffArea 0.373 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.485 1.750 4.735 1.930 ;
        RECT  4.365 1.750 4.485 2.140 ;
        RECT  3.235 2.020 4.365 2.140 ;
        RECT  3.065 2.020 3.235 2.190 ;
        END
        AntennaGateArea 0.1814 ;
    END CS
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 0.450 0.590 0.710 ;
        RECT  0.375 0.450 0.490 0.775 ;
        RECT  0.195 0.655 0.375 0.775 ;
        RECT  0.195 1.425 0.230 2.045 ;
        RECT  0.070 0.655 0.195 2.045 ;
        END
        AntennaDiffArea 0.354 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.530 1.900 2.940 2.020 ;
        RECT  1.410 0.980 1.530 2.020 ;
        RECT  1.350 0.980 1.410 1.240 ;
        RECT  0.490 1.735 1.410 1.855 ;
        RECT  0.350 1.010 0.490 1.855 ;
        RECT  0.320 1.010 0.350 1.270 ;
        END
        AntennaGateArea 0.3508 ;
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.050 1.200 1.235 ;
        RECT  0.910 1.050 1.050 1.375 ;
        END
        AntennaGateArea 0.1629 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.850 -0.210 5.320 0.210 ;
        RECT  4.590 -0.210 4.850 0.230 ;
        RECT  2.630 -0.210 4.590 0.210 ;
        RECT  2.370 -0.210 2.630 0.320 ;
        RECT  1.020 -0.210 2.370 0.210 ;
        RECT  0.760 -0.210 1.020 0.500 ;
        RECT  0.255 -0.210 0.760 0.210 ;
        RECT  0.085 -0.210 0.255 0.535 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.875 2.310 5.320 2.730 ;
        RECT  4.705 2.105 4.875 2.730 ;
        RECT  2.680 2.310 4.705 2.730 ;
        RECT  2.420 2.140 2.680 2.730 ;
        RECT  0.915 2.310 2.420 2.730 ;
        RECT  0.745 1.975 0.915 2.730 ;
        RECT  0.000 2.310 0.745 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.320 2.520 ;
        LAYER M1 ;
        RECT  4.850 0.380 4.970 1.270 ;
        RECT  3.685 0.380 4.850 0.500 ;
        RECT  4.485 0.620 4.530 0.740 ;
        RECT  4.315 0.620 4.485 1.600 ;
        RECT  4.270 0.620 4.315 0.740 ;
        RECT  4.220 1.070 4.315 1.330 ;
        RECT  4.070 1.730 4.145 1.900 ;
        RECT  4.070 0.620 4.115 0.740 ;
        RECT  3.950 0.620 4.070 1.900 ;
        RECT  3.855 0.620 3.950 0.740 ;
        RECT  3.245 1.780 3.950 1.900 ;
        RECT  3.685 1.540 3.830 1.660 ;
        RECT  3.565 0.380 3.685 1.660 ;
        RECT  3.320 1.420 3.400 1.540 ;
        RECT  3.200 0.440 3.320 1.540 ;
        RECT  3.125 1.660 3.245 1.900 ;
        RECT  2.250 0.440 3.200 0.560 ;
        RECT  3.140 1.420 3.200 1.540 ;
        RECT  1.770 1.660 3.125 1.780 ;
        RECT  2.870 1.325 3.015 1.495 ;
        RECT  2.870 0.680 3.010 0.800 ;
        RECT  2.750 0.680 2.870 1.495 ;
        RECT  2.010 1.375 2.750 1.495 ;
        RECT  2.250 0.960 2.340 1.220 ;
        RECT  2.130 0.440 2.250 1.220 ;
        RECT  2.040 0.440 2.130 0.560 ;
        RECT  1.905 0.380 2.040 0.560 ;
        RECT  1.890 0.980 2.010 1.495 ;
        RECT  1.365 0.380 1.905 0.500 ;
        RECT  1.650 0.625 1.770 1.780 ;
        RECT  1.600 0.625 1.650 0.795 ;
        RECT  1.195 0.380 1.365 0.740 ;
        RECT  1.170 1.355 1.290 1.615 ;
        RECT  0.830 0.620 1.195 0.740 ;
        RECT  0.770 1.495 1.170 1.615 ;
        RECT  0.770 0.620 0.830 0.945 ;
        RECT  0.710 0.620 0.770 1.615 ;
        RECT  0.650 0.825 0.710 1.615 ;
    END
END AHCSHCINX2AD
MACRO AHCSHCINX4AD
    CLASS CORE ;
    FOREIGN AHCSHCINX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.930 0.400 6.090 1.965 ;
        END
        AntennaDiffArea 0.373 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.135 1.750 5.400 1.930 ;
        RECT  5.015 1.750 5.135 2.140 ;
        RECT  3.945 2.020 5.015 2.140 ;
        RECT  3.775 2.020 3.945 2.190 ;
        END
        AntennaGateArea 0.181 ;
    END CS
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.385 1.310 0.645 ;
        RECT  0.515 0.525 1.190 0.645 ;
        RECT  0.805 1.420 0.975 2.065 ;
        RECT  0.210 1.420 0.805 1.560 ;
        RECT  0.375 0.525 0.515 0.865 ;
        RECT  0.210 0.725 0.375 0.865 ;
        RECT  0.070 0.725 0.210 1.560 ;
        END
        AntennaDiffArea 0.522 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.180 1.900 3.650 2.020 ;
        RECT  2.060 0.980 2.180 2.020 ;
        RECT  1.655 1.770 2.060 1.895 ;
        RECT  1.220 1.750 1.655 1.895 ;
        RECT  1.100 1.080 1.220 1.895 ;
        RECT  0.875 1.080 1.100 1.250 ;
        END
        AntennaGateArea 0.4978 ;
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.865 1.890 1.270 ;
        RECT  1.630 1.080 1.750 1.270 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 -0.210 6.160 0.210 ;
        RECT  5.570 -0.210 5.690 0.720 ;
        RECT  3.340 -0.210 5.570 0.210 ;
        RECT  3.080 -0.210 3.340 0.320 ;
        RECT  1.740 -0.210 3.080 0.210 ;
        RECT  1.480 -0.210 1.740 0.390 ;
        RECT  1.020 -0.210 1.480 0.210 ;
        RECT  0.760 -0.210 1.020 0.390 ;
        RECT  0.255 -0.210 0.760 0.210 ;
        RECT  0.085 -0.210 0.255 0.605 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 2.310 6.160 2.730 ;
        RECT  5.545 1.585 5.715 2.730 ;
        RECT  3.390 2.310 5.545 2.730 ;
        RECT  3.130 2.140 3.390 2.730 ;
        RECT  1.630 2.310 3.130 2.730 ;
        RECT  1.370 2.025 1.630 2.730 ;
        RECT  0.365 2.310 1.370 2.730 ;
        RECT  0.195 1.690 0.365 2.730 ;
        RECT  0.000 2.310 0.195 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.690 1.010 5.810 1.270 ;
        RECT  5.450 1.010 5.690 1.130 ;
        RECT  5.330 0.380 5.450 1.130 ;
        RECT  4.400 0.380 5.330 0.500 ;
        RECT  5.040 0.620 5.210 1.600 ;
        RECT  4.950 0.620 5.040 0.740 ;
        RECT  4.975 1.070 5.040 1.330 ;
        RECT  4.710 0.620 4.830 1.900 ;
        RECT  4.570 0.620 4.710 0.740 ;
        RECT  3.890 1.780 4.710 1.900 ;
        RECT  4.400 1.540 4.540 1.660 ;
        RECT  4.280 0.380 4.400 1.660 ;
        RECT  4.035 1.420 4.110 1.540 ;
        RECT  3.915 0.440 4.035 1.540 ;
        RECT  3.050 0.440 3.915 0.560 ;
        RECT  3.850 1.420 3.915 1.540 ;
        RECT  3.770 1.660 3.890 1.900 ;
        RECT  2.480 1.660 3.770 1.780 ;
        RECT  3.580 1.325 3.725 1.495 ;
        RECT  3.580 0.680 3.720 0.800 ;
        RECT  3.460 0.680 3.580 1.495 ;
        RECT  2.720 1.375 3.460 1.495 ;
        RECT  2.930 0.440 3.050 1.220 ;
        RECT  2.800 0.440 2.930 0.560 ;
        RECT  2.620 0.380 2.800 0.560 ;
        RECT  2.600 0.980 2.720 1.495 ;
        RECT  2.055 0.380 2.620 0.500 ;
        RECT  2.360 0.625 2.480 1.780 ;
        RECT  2.310 0.625 2.360 0.795 ;
        RECT  1.885 0.380 2.055 0.745 ;
        RECT  1.810 1.390 1.940 1.650 ;
        RECT  1.550 0.625 1.885 0.745 ;
        RECT  1.460 1.390 1.810 1.510 ;
        RECT  1.460 0.625 1.550 0.890 ;
        RECT  1.430 0.625 1.460 1.510 ;
        RECT  1.340 0.770 1.430 1.510 ;
        RECT  0.755 0.770 1.340 0.890 ;
        RECT  0.635 0.770 0.755 1.160 ;
        RECT  0.450 1.040 0.635 1.160 ;
        RECT  0.330 1.040 0.450 1.300 ;
    END
END AHCSHCINX4AD
MACRO AHCSHCONX2AD
    CLASS CORE ;
    FOREIGN AHCSHCONX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.090 0.400 5.250 1.965 ;
        END
        AntennaDiffArea 0.373 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.355 1.750 4.735 1.930 ;
        RECT  4.235 1.750 4.355 2.140 ;
        RECT  3.015 2.020 4.235 2.140 ;
        END
        AntennaGateArea 0.1814 ;
    END CS
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.445 1.600 0.615 2.055 ;
        RECT  0.210 1.600 0.445 1.720 ;
        RECT  0.210 0.415 0.290 0.845 ;
        RECT  0.120 0.415 0.210 1.720 ;
        RECT  0.070 0.650 0.120 1.720 ;
        END
        AntennaDiffArea 0.343 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.935 2.020 2.895 2.140 ;
        RECT  1.705 2.020 1.935 2.170 ;
        RECT  1.550 2.020 1.705 2.140 ;
        RECT  1.430 1.140 1.550 2.140 ;
        RECT  0.895 1.820 1.430 1.940 ;
        RECT  0.775 1.360 0.895 1.940 ;
        RECT  0.450 1.360 0.775 1.480 ;
        RECT  0.330 1.030 0.450 1.480 ;
        END
        AntennaGateArea 0.3399 ;
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.980 1.200 ;
        END
        AntennaGateArea 0.302 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.850 -0.210 5.320 0.210 ;
        RECT  4.590 -0.210 4.850 0.230 ;
        RECT  2.670 -0.210 4.590 0.210 ;
        RECT  2.410 -0.210 2.670 0.380 ;
        RECT  0.935 -0.210 2.410 0.210 ;
        RECT  0.765 -0.210 0.935 0.710 ;
        RECT  0.000 -0.210 0.765 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.875 2.310 5.320 2.730 ;
        RECT  4.705 2.105 4.875 2.730 ;
        RECT  2.590 2.310 4.705 2.730 ;
        RECT  2.420 2.265 2.590 2.730 ;
        RECT  1.020 2.310 2.420 2.730 ;
        RECT  0.760 2.070 1.020 2.730 ;
        RECT  0.255 2.310 0.760 2.730 ;
        RECT  0.085 1.840 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.320 2.520 ;
        LAYER M1 ;
        RECT  4.850 0.380 4.970 1.270 ;
        RECT  3.680 0.380 4.850 0.500 ;
        RECT  4.480 0.620 4.525 0.740 ;
        RECT  4.310 0.620 4.480 1.600 ;
        RECT  4.265 0.620 4.310 0.740 ;
        RECT  4.185 1.070 4.310 1.330 ;
        RECT  4.065 1.640 4.115 1.900 ;
        RECT  4.065 0.620 4.110 0.740 ;
        RECT  3.945 0.620 4.065 1.900 ;
        RECT  3.850 0.620 3.945 0.740 ;
        RECT  1.790 1.780 3.945 1.900 ;
        RECT  3.680 1.540 3.825 1.660 ;
        RECT  3.560 0.380 3.680 1.660 ;
        RECT  3.320 1.540 3.440 1.660 ;
        RECT  3.180 0.500 3.320 1.660 ;
        RECT  2.370 0.500 3.180 0.620 ;
        RECT  2.930 0.740 3.050 1.660 ;
        RECT  2.790 0.740 2.930 0.860 ;
        RECT  2.035 1.540 2.930 1.660 ;
        RECT  2.250 0.500 2.370 1.395 ;
        RECT  2.125 0.500 2.250 0.620 ;
        RECT  2.005 0.380 2.125 0.620 ;
        RECT  1.915 1.190 2.035 1.660 ;
        RECT  1.335 0.380 2.005 0.500 ;
        RECT  1.790 0.645 1.840 0.815 ;
        RECT  1.670 0.645 1.790 1.900 ;
        RECT  1.285 0.380 1.335 0.810 ;
        RECT  1.285 1.400 1.310 1.660 ;
        RECT  1.165 0.380 1.285 1.660 ;
    END
END AHCSHCONX2AD
MACRO AHCSHCONX4AD
    CLASS CORE ;
    FOREIGN AHCSHCONX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.930 0.400 6.090 1.965 ;
        END
        AntennaDiffArea 0.373 ;
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.145 1.750 5.575 1.930 ;
        RECT  5.025 1.750 5.145 2.140 ;
        RECT  3.805 2.020 5.025 2.140 ;
        END
        AntennaGateArea 0.1814 ;
    END CS
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.165 1.600 1.335 2.030 ;
        RECT  0.615 1.600 1.165 1.730 ;
        RECT  0.815 0.550 0.985 0.750 ;
        RECT  0.210 0.620 0.815 0.750 ;
        RECT  0.445 1.600 0.615 2.030 ;
        RECT  0.210 1.600 0.445 1.730 ;
        RECT  0.070 0.620 0.210 1.730 ;
        END
        AntennaDiffArea 0.562 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.775 2.020 3.685 2.140 ;
        RECT  2.545 2.020 2.775 2.170 ;
        RECT  2.340 2.020 2.545 2.140 ;
        RECT  2.220 1.140 2.340 2.140 ;
        RECT  1.620 1.775 2.220 1.900 ;
        RECT  1.500 1.360 1.620 1.900 ;
        RECT  1.130 1.360 1.500 1.480 ;
        RECT  0.910 1.110 1.130 1.480 ;
        RECT  0.610 1.110 0.910 1.255 ;
        END
        AntennaGateArea 0.4799 ;
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.395 0.630 1.655 1.230 ;
        RECT  0.450 0.870 1.395 0.990 ;
        RECT  0.330 0.870 0.450 1.280 ;
        END
        AntennaGateArea 0.442 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.690 -0.210 6.160 0.210 ;
        RECT  5.430 -0.210 5.690 0.230 ;
        RECT  3.460 -0.210 5.430 0.210 ;
        RECT  3.200 -0.210 3.460 0.380 ;
        RECT  1.655 -0.210 3.200 0.210 ;
        RECT  1.395 -0.210 1.655 0.510 ;
        RECT  0.410 -0.210 1.395 0.210 ;
        RECT  0.150 -0.210 0.410 0.500 ;
        RECT  0.000 -0.210 0.150 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.665 2.310 6.160 2.730 ;
        RECT  5.495 2.105 5.665 2.730 ;
        RECT  3.380 2.310 5.495 2.730 ;
        RECT  3.210 2.265 3.380 2.730 ;
        RECT  1.740 2.310 3.210 2.730 ;
        RECT  1.480 2.020 1.740 2.730 ;
        RECT  0.975 2.310 1.480 2.730 ;
        RECT  0.805 1.850 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.850 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.690 0.380 5.810 1.270 ;
        RECT  4.470 0.380 5.690 0.500 ;
        RECT  5.270 0.620 5.315 0.740 ;
        RECT  5.100 0.620 5.270 1.600 ;
        RECT  5.055 0.620 5.100 0.740 ;
        RECT  4.975 1.070 5.100 1.330 ;
        RECT  4.855 1.640 4.905 1.900 ;
        RECT  4.855 0.620 4.900 0.740 ;
        RECT  4.735 0.620 4.855 1.900 ;
        RECT  4.640 0.620 4.735 0.740 ;
        RECT  2.580 1.780 4.735 1.900 ;
        RECT  4.470 1.540 4.615 1.660 ;
        RECT  4.350 0.380 4.470 1.660 ;
        RECT  4.110 1.540 4.230 1.660 ;
        RECT  3.990 0.500 4.110 1.660 ;
        RECT  3.195 0.500 3.990 0.620 ;
        RECT  3.970 1.540 3.990 1.660 ;
        RECT  3.720 0.740 3.840 1.660 ;
        RECT  3.580 0.740 3.720 0.860 ;
        RECT  2.825 1.540 3.720 1.660 ;
        RECT  3.160 0.500 3.195 1.305 ;
        RECT  3.075 0.500 3.160 1.395 ;
        RECT  2.885 0.500 3.075 0.620 ;
        RECT  3.040 1.135 3.075 1.395 ;
        RECT  2.765 0.380 2.885 0.620 ;
        RECT  2.705 1.190 2.825 1.660 ;
        RECT  2.010 0.380 2.765 0.500 ;
        RECT  2.580 0.645 2.630 0.815 ;
        RECT  2.460 0.645 2.580 1.900 ;
        RECT  2.010 1.535 2.100 1.655 ;
        RECT  1.890 0.380 2.010 1.655 ;
        RECT  1.840 1.535 1.890 1.655 ;
    END
END AHCSHCONX4AD
MACRO AHHCINX2AD
    CLASS CORE ;
    FOREIGN AHHCINX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.145 2.170 1.750 ;
        RECT  1.980 0.665 2.120 1.750 ;
        RECT  1.860 0.665 1.980 0.925 ;
        RECT  1.930 1.510 1.980 1.750 ;
        RECT  1.350 1.510 1.930 1.630 ;
        RECT  1.180 1.460 1.350 1.630 ;
        END
        AntennaDiffArea 0.536 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.045 0.700 4.130 1.740 ;
        RECT  3.990 0.700 4.045 2.010 ;
        RECT  3.840 0.700 3.990 0.820 ;
        RECT  3.875 1.580 3.990 2.010 ;
        RECT  3.720 0.515 3.840 0.820 ;
        RECT  3.540 0.515 3.720 0.635 ;
        END
        AntennaDiffArea 0.392 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.405 1.425 3.570 2.020 ;
        RECT  3.360 1.235 3.405 2.020 ;
        RECT  3.285 1.030 3.360 2.020 ;
        RECT  3.240 1.030 3.285 1.355 ;
        RECT  2.095 1.900 3.285 2.020 ;
        RECT  1.975 1.900 2.095 2.140 ;
        RECT  1.125 2.020 1.975 2.140 ;
        RECT  0.955 2.020 1.125 2.190 ;
        END
        AntennaGateArea 0.3835 ;
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.865 2.730 1.375 ;
        END
        AntennaGateArea 0.2327 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.100 -0.210 4.200 0.210 ;
        RECT  3.960 -0.210 4.100 0.580 ;
        RECT  3.205 -0.210 3.960 0.210 ;
        RECT  2.775 -0.210 3.205 0.365 ;
        RECT  0.730 -0.210 2.775 0.210 ;
        RECT  0.470 -0.210 0.730 0.310 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.365 2.310 4.200 2.730 ;
        RECT  3.195 2.190 3.365 2.730 ;
        RECT  2.840 2.310 3.195 2.730 ;
        RECT  2.670 2.190 2.840 2.730 ;
        RECT  0.660 2.310 2.670 2.730 ;
        RECT  0.540 2.150 0.660 2.730 ;
        RECT  0.000 2.310 0.540 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  3.750 0.940 3.870 1.280 ;
        RECT  3.600 0.940 3.750 1.060 ;
        RECT  3.480 0.755 3.600 1.060 ;
        RECT  3.090 0.755 3.480 0.875 ;
        RECT  3.090 1.505 3.125 1.765 ;
        RECT  2.970 0.680 3.090 1.765 ;
        RECT  2.930 0.680 2.970 0.940 ;
        RECT  2.340 0.420 2.460 1.720 ;
        RECT  2.240 0.420 2.340 0.940 ;
        RECT  2.290 1.550 2.340 1.720 ;
        RECT  1.740 0.420 2.240 0.540 ;
        RECT  0.255 1.780 1.785 1.900 ;
        RECT  1.505 1.170 1.765 1.380 ;
        RECT  1.620 0.420 1.740 1.050 ;
        RECT  0.680 0.930 1.620 1.050 ;
        RECT  1.045 1.170 1.505 1.290 ;
        RECT  1.380 0.430 1.500 0.755 ;
        RECT  0.255 0.430 1.380 0.550 ;
        RECT  0.440 0.680 1.230 0.800 ;
        RECT  0.925 1.170 1.045 1.660 ;
        RECT  0.785 1.420 0.925 1.660 ;
        RECT  0.440 1.420 0.785 1.540 ;
        RECT  0.560 0.930 0.680 1.210 ;
        RECT  0.320 0.680 0.440 1.540 ;
        RECT  0.200 0.380 0.255 0.550 ;
        RECT  0.200 1.780 0.255 1.950 ;
        RECT  0.080 0.380 0.200 1.950 ;
    END
END AHHCINX2AD
MACRO AHHCINX4AD
    CLASS CORE ;
    FOREIGN AHHCINX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.005 2.170 1.750 ;
        RECT  1.980 0.665 2.120 1.750 ;
        RECT  1.860 0.665 1.980 0.925 ;
        RECT  1.930 1.510 1.980 1.750 ;
        RECT  1.350 1.510 1.930 1.630 ;
        RECT  1.180 1.460 1.350 1.630 ;
        END
        AntennaDiffArea 0.536 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.830 0.540 4.970 1.740 ;
        RECT  4.625 0.540 4.830 0.680 ;
        RECT  4.210 1.580 4.830 1.740 ;
        RECT  4.365 0.510 4.625 0.680 ;
        RECT  3.625 0.510 4.365 0.650 ;
        RECT  4.040 1.580 4.210 2.010 ;
        END
        AntennaDiffArea 0.618 ;
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.525 1.015 4.665 1.455 ;
        RECT  3.665 1.315 4.525 1.455 ;
        RECT  3.570 1.010 3.665 1.455 ;
        RECT  3.410 1.010 3.570 2.020 ;
        RECT  2.095 1.900 3.410 2.020 ;
        RECT  1.975 1.900 2.095 2.140 ;
        RECT  1.125 2.020 1.975 2.140 ;
        RECT  0.955 2.020 1.125 2.190 ;
        END
        AntennaGateArea 0.5445 ;
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.865 2.730 1.375 ;
        END
        AntennaGateArea 0.3091 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.940 -0.210 5.040 0.210 ;
        RECT  4.770 -0.210 4.940 0.415 ;
        RECT  4.245 -0.210 4.770 0.210 ;
        RECT  3.985 -0.210 4.245 0.390 ;
        RECT  3.480 -0.210 3.985 0.210 ;
        RECT  3.310 -0.210 3.480 0.415 ;
        RECT  2.815 -0.210 3.310 0.210 ;
        RECT  2.645 -0.210 2.815 0.365 ;
        RECT  0.730 -0.210 2.645 0.210 ;
        RECT  0.470 -0.210 0.730 0.310 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.875 2.310 5.040 2.730 ;
        RECT  4.615 1.870 4.875 2.730 ;
        RECT  3.505 2.310 4.615 2.730 ;
        RECT  3.335 2.190 3.505 2.730 ;
        RECT  2.840 2.310 3.335 2.730 ;
        RECT  2.670 2.190 2.840 2.730 ;
        RECT  0.660 2.310 2.670 2.730 ;
        RECT  0.540 2.150 0.660 2.730 ;
        RECT  0.000 2.310 0.540 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.040 2.520 ;
        LAYER M1 ;
        RECT  4.000 1.025 4.340 1.195 ;
        RECT  3.880 0.770 4.000 1.195 ;
        RECT  3.170 0.770 3.880 0.890 ;
        RECT  3.090 1.505 3.195 1.765 ;
        RECT  3.090 0.680 3.170 0.940 ;
        RECT  2.970 0.680 3.090 1.765 ;
        RECT  2.340 0.420 2.460 1.720 ;
        RECT  2.240 0.420 2.340 0.770 ;
        RECT  2.290 1.550 2.340 1.720 ;
        RECT  1.740 0.420 2.240 0.540 ;
        RECT  0.255 1.780 1.785 1.900 ;
        RECT  1.505 1.170 1.765 1.380 ;
        RECT  1.620 0.420 1.740 1.050 ;
        RECT  0.680 0.930 1.620 1.050 ;
        RECT  1.045 1.170 1.505 1.290 ;
        RECT  1.380 0.430 1.500 0.755 ;
        RECT  0.255 0.430 1.380 0.550 ;
        RECT  0.440 0.680 1.230 0.800 ;
        RECT  0.925 1.170 1.045 1.660 ;
        RECT  0.785 1.420 0.925 1.660 ;
        RECT  0.440 1.420 0.785 1.540 ;
        RECT  0.560 0.930 0.680 1.210 ;
        RECT  0.320 0.680 0.440 1.540 ;
        RECT  0.200 0.380 0.255 0.550 ;
        RECT  0.200 1.780 0.255 1.950 ;
        RECT  0.080 0.380 0.200 1.950 ;
    END
END AHHCINX4AD
MACRO AHHCONX2AD
    CLASS CORE ;
    FOREIGN AHHCONX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.835 1.775 1.925 1.895 ;
        RECT  1.715 0.620 1.835 1.895 ;
        RECT  1.665 1.425 1.715 1.895 ;
        RECT  1.470 1.425 1.665 1.655 ;
        END
        AntennaDiffArea 0.516 ;
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.760 3.570 1.735 ;
        RECT  3.430 0.405 3.450 1.735 ;
        RECT  3.280 0.405 3.430 0.880 ;
        RECT  3.195 1.615 3.430 1.735 ;
        RECT  3.025 1.615 3.195 2.045 ;
        END
        AntennaDiffArea 0.443 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.000 3.295 1.410 ;
        RECT  2.560 1.290 3.150 1.410 ;
        RECT  2.440 1.290 2.560 1.985 ;
        RECT  2.315 1.290 2.440 1.410 ;
        RECT  2.320 1.865 2.440 2.140 ;
        RECT  0.730 2.020 2.320 2.140 ;
        RECT  2.195 1.005 2.315 1.410 ;
        END
        AntennaGateArea 0.358 ;
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.865 2.975 1.170 ;
        RECT  2.455 1.050 2.590 1.170 ;
        END
        AntennaGateArea 0.324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.885 -0.210 3.640 0.210 ;
        RECT  2.625 -0.210 2.885 0.715 ;
        RECT  0.750 -0.210 2.625 0.210 ;
        RECT  0.490 -0.210 0.750 0.310 ;
        RECT  0.000 -0.210 0.490 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.555 2.310 3.640 2.730 ;
        RECT  3.385 1.855 3.555 2.730 ;
        RECT  2.790 2.310 3.385 2.730 ;
        RECT  2.620 2.105 2.790 2.730 ;
        RECT  0.610 2.310 2.620 2.730 ;
        RECT  0.420 2.020 0.610 2.730 ;
        RECT  0.000 2.310 0.420 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  2.075 0.470 2.480 0.640 ;
        RECT  2.150 1.535 2.320 1.705 ;
        RECT  2.075 1.535 2.150 1.655 ;
        RECT  1.955 0.380 2.075 1.655 ;
        RECT  1.575 0.380 1.955 0.500 ;
        RECT  1.455 0.380 1.575 1.040 ;
        RECT  0.275 1.780 1.545 1.900 ;
        RECT  0.710 0.920 1.455 1.040 ;
        RECT  1.285 1.160 1.445 1.280 ;
        RECT  1.075 0.340 1.335 0.560 ;
        RECT  1.230 1.160 1.285 1.520 ;
        RECT  0.470 0.680 1.230 0.800 ;
        RECT  1.165 1.160 1.230 1.560 ;
        RECT  0.970 1.400 1.165 1.560 ;
        RECT  0.275 0.440 1.075 0.560 ;
        RECT  0.470 1.400 0.970 1.520 ;
        RECT  0.590 0.920 0.710 1.270 ;
        RECT  0.350 0.680 0.470 1.520 ;
        RECT  0.230 0.390 0.275 0.560 ;
        RECT  0.230 1.725 0.275 2.155 ;
        RECT  0.105 0.390 0.230 2.155 ;
    END
END AHHCONX2AD
MACRO AHHCONX4AD
    CLASS CORE ;
    FOREIGN AHHCONX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.115 0.630 3.255 1.220 ;
        RECT  3.070 1.640 3.190 1.900 ;
        RECT  2.470 1.060 3.115 1.220 ;
        RECT  2.470 1.775 3.070 1.900 ;
        RECT  2.450 1.060 2.470 1.900 ;
        RECT  2.310 0.860 2.450 1.900 ;
        RECT  1.950 0.860 2.310 1.000 ;
        RECT  1.560 1.500 2.310 1.640 ;
        END
        AntennaDiffArea 0.928 ;
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.955 0.625 6.090 1.685 ;
        RECT  5.950 0.345 5.955 1.685 ;
        RECT  5.835 0.345 5.950 0.865 ;
        RECT  5.675 1.545 5.950 1.685 ;
        RECT  4.745 0.625 5.835 0.765 ;
        RECT  5.505 1.545 5.675 1.995 ;
        RECT  4.880 1.545 5.505 1.685 ;
        RECT  4.710 1.545 4.880 1.995 ;
        RECT  4.485 0.385 4.745 0.765 ;
        END
        AntennaDiffArea 0.952 ;
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.685 1.020 5.805 1.425 ;
        RECT  4.890 1.305 5.685 1.425 ;
        RECT  4.505 1.125 4.890 1.425 ;
        RECT  4.380 1.305 4.505 1.425 ;
        RECT  4.260 1.305 4.380 1.760 ;
        RECT  3.450 1.640 4.260 1.760 ;
        RECT  3.330 1.640 3.450 2.170 ;
        RECT  1.630 2.020 3.330 2.140 ;
        RECT  1.370 2.020 1.630 2.190 ;
        END
        AntennaGateArea 0.7092 ;
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.245 1.065 5.535 1.185 ;
        RECT  5.015 0.885 5.245 1.185 ;
        RECT  4.180 0.885 5.015 1.005 ;
        RECT  3.750 0.885 4.180 1.210 ;
        END
        AntennaGateArea 0.648 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.385 -0.210 6.160 0.210 ;
        RECT  5.125 -0.210 5.385 0.505 ;
        RECT  4.035 -0.210 5.125 0.210 ;
        RECT  3.775 -0.210 4.035 0.525 ;
        RECT  1.040 -0.210 3.775 0.210 ;
        RECT  0.780 -0.210 1.040 0.310 ;
        RECT  0.230 -0.210 0.780 0.210 ;
        RECT  0.110 -0.210 0.230 0.885 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.040 2.310 6.160 2.730 ;
        RECT  5.870 1.805 6.040 2.730 ;
        RECT  5.310 2.310 5.870 2.730 ;
        RECT  5.140 1.805 5.310 2.730 ;
        RECT  4.455 2.310 5.140 2.730 ;
        RECT  4.285 1.880 4.455 2.730 ;
        RECT  3.735 2.310 4.285 2.730 ;
        RECT  3.570 1.880 3.735 2.730 ;
        RECT  1.050 2.310 3.570 2.730 ;
        RECT  0.790 2.210 1.050 2.730 ;
        RECT  0.230 2.310 0.790 2.730 ;
        RECT  0.110 1.520 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  4.180 0.595 4.350 0.765 ;
        RECT  3.630 0.645 4.180 0.765 ;
        RECT  3.630 1.400 4.140 1.520 ;
        RECT  3.460 0.380 3.630 1.520 ;
        RECT  2.885 0.380 3.460 0.500 ;
        RECT  2.900 1.400 3.460 1.520 ;
        RECT  2.640 1.400 2.900 1.655 ;
        RECT  2.765 0.380 2.885 0.740 ;
        RECT  1.710 0.620 2.765 0.740 ;
        RECT  1.345 0.380 2.600 0.500 ;
        RECT  0.470 1.780 2.180 1.900 ;
        RECT  1.590 0.620 1.710 1.040 ;
        RECT  1.400 1.160 1.700 1.280 ;
        RECT  0.950 0.920 1.590 1.040 ;
        RECT  0.710 0.680 1.470 0.800 ;
        RECT  1.280 1.160 1.400 1.645 ;
        RECT  1.205 0.380 1.345 0.550 ;
        RECT  0.710 1.525 1.280 1.645 ;
        RECT  0.470 0.430 1.205 0.550 ;
        RECT  0.830 0.920 0.950 1.260 ;
        RECT  0.590 0.680 0.710 1.645 ;
        RECT  0.350 0.430 0.470 1.900 ;
    END
END AHHCONX4AD
MACRO AND2X1AD
    CLASS CORE ;
    FOREIGN AND2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.640 1.330 1.935 ;
        END
        AntennaDiffArea 0.216 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.020 0.770 1.375 ;
        END
        AntennaGateArea 0.0424 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.055 0.365 1.315 ;
        RECT  0.070 1.055 0.210 1.655 ;
        END
        AntennaGateArea 0.0424 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 -0.210 1.400 0.210 ;
        RECT  0.750 -0.210 0.920 0.660 ;
        RECT  0.000 -0.210 0.750 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.925 2.310 1.400 2.730 ;
        RECT  0.755 1.925 0.925 2.730 ;
        RECT  0.255 2.310 0.755 2.730 ;
        RECT  0.085 1.925 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.920 0.780 1.040 1.615 ;
        RECT  0.270 0.780 0.920 0.900 ;
        RECT  0.390 1.495 0.920 1.615 ;
        RECT  0.100 0.730 0.270 0.900 ;
    END
END AND2X1AD
MACRO AND2X2AD
    CLASS CORE ;
    FOREIGN AND2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.430 1.330 1.935 ;
        END
        AntennaDiffArea 0.389 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.020 0.770 1.375 ;
        END
        AntennaGateArea 0.0754 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.065 0.320 1.235 ;
        RECT  0.070 1.065 0.210 1.655 ;
        END
        AntennaGateArea 0.0754 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.965 -0.210 1.400 0.210 ;
        RECT  0.705 -0.210 0.965 0.650 ;
        RECT  0.000 -0.210 0.705 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.925 2.310 1.400 2.730 ;
        RECT  0.755 1.985 0.925 2.730 ;
        RECT  0.255 2.310 0.755 2.730 ;
        RECT  0.085 1.985 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.920 0.780 1.040 1.615 ;
        RECT  0.270 0.780 0.920 0.900 ;
        RECT  0.390 1.495 0.920 1.615 ;
        RECT  0.100 0.730 0.270 0.900 ;
    END
END AND2X2AD
MACRO AND2X4AD
    CLASS CORE ;
    FOREIGN AND2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 1.005 1.890 1.515 ;
        RECT  1.640 0.420 1.760 2.060 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.280 1.250 1.400 ;
        RECT  0.210 1.140 0.330 1.400 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.147 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.780 0.910 1.095 1.050 ;
        RECT  0.520 0.910 0.780 1.160 ;
        END
        AntennaGateArea 0.147 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.120 -0.210 2.240 0.210 ;
        RECT  2.000 -0.210 2.120 0.830 ;
        RECT  1.355 -0.210 2.000 0.210 ;
        RECT  1.185 -0.210 1.355 0.315 ;
        RECT  0.260 -0.210 1.185 0.210 ;
        RECT  0.090 -0.210 0.260 0.315 ;
        RECT  0.000 -0.210 0.090 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.120 2.310 2.240 2.730 ;
        RECT  2.000 1.690 2.120 2.730 ;
        RECT  1.470 2.310 2.000 2.730 ;
        RECT  1.210 1.870 1.470 2.730 ;
        RECT  1.020 2.310 1.210 2.730 ;
        RECT  0.760 1.870 1.020 2.730 ;
        RECT  0.230 2.310 0.760 2.730 ;
        RECT  0.110 1.770 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.400 0.650 1.520 1.740 ;
        RECT  0.620 0.650 1.400 0.770 ;
        RECT  0.615 1.620 1.400 1.740 ;
        RECT  0.445 1.620 0.615 2.050 ;
    END
END AND2X4AD
MACRO AND2X6AD
    CLASS CORE ;
    FOREIGN AND2X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 0.345 2.730 2.030 ;
        RECT  2.560 0.670 2.570 1.565 ;
        RECT  1.995 0.670 2.560 0.865 ;
        RECT  1.995 1.385 2.560 1.565 ;
        RECT  1.825 0.435 1.995 0.865 ;
        RECT  1.825 1.385 1.995 1.990 ;
        END
        AntennaDiffArea 0.795 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.235 1.020 1.355 1.410 ;
        RECT  0.210 1.290 1.235 1.410 ;
        RECT  0.070 1.020 0.210 1.655 ;
        END
        AntennaGateArea 0.2229 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.575 0.910 1.095 1.170 ;
        END
        AntennaGateArea 0.2228 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.400 -0.210 2.800 0.210 ;
        RECT  2.140 -0.210 2.400 0.500 ;
        RECT  1.615 -0.210 2.140 0.210 ;
        RECT  1.445 -0.210 1.615 0.555 ;
        RECT  0.255 -0.210 1.445 0.210 ;
        RECT  0.085 -0.210 0.255 0.815 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.355 2.310 2.800 2.730 ;
        RECT  2.185 1.840 2.355 2.730 ;
        RECT  1.565 2.310 2.185 2.730 ;
        RECT  1.395 2.165 1.565 2.730 ;
        RECT  0.935 2.310 1.395 2.730 ;
        RECT  0.765 2.165 0.935 2.730 ;
        RECT  0.255 2.310 0.765 2.730 ;
        RECT  0.085 2.165 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  1.595 1.040 2.195 1.185 ;
        RECT  1.475 0.715 1.595 1.700 ;
        RECT  1.325 0.715 1.475 0.835 ;
        RECT  0.430 1.530 1.475 1.700 ;
        RECT  1.205 0.620 1.325 0.835 ;
        RECT  0.910 0.620 1.205 0.740 ;
        RECT  0.740 0.555 0.910 0.740 ;
    END
END AND2X6AD
MACRO AND2X8AD
    CLASS CORE ;
    FOREIGN AND2X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 0.620 3.710 1.590 ;
        RECT  3.260 0.420 3.430 1.960 ;
        RECT  2.710 0.620 3.260 0.870 ;
        RECT  2.710 1.340 3.260 1.590 ;
        RECT  2.540 0.420 2.710 0.870 ;
        RECT  2.535 1.340 2.710 1.965 ;
        END
        AntennaDiffArea 0.844 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.185 1.290 2.105 1.410 ;
        RECT  0.865 1.110 1.185 1.410 ;
        RECT  0.665 1.110 0.865 1.230 ;
        END
        AntennaGateArea 0.2948 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.455 1.040 1.590 1.160 ;
        RECT  1.330 0.865 1.455 1.160 ;
        RECT  0.490 0.865 1.330 0.990 ;
        RECT  0.335 0.865 0.490 1.375 ;
        END
        AntennaGateArea 0.294 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.790 -0.210 3.920 0.210 ;
        RECT  3.620 -0.210 3.790 0.500 ;
        RECT  3.115 -0.210 3.620 0.210 ;
        RECT  2.855 -0.210 3.115 0.500 ;
        RECT  2.350 -0.210 2.855 0.210 ;
        RECT  2.180 -0.210 2.350 0.675 ;
        RECT  1.070 -0.210 2.180 0.210 ;
        RECT  0.810 -0.210 1.070 0.505 ;
        RECT  0.000 -0.210 0.810 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.790 2.310 3.920 2.730 ;
        RECT  3.620 1.845 3.790 2.730 ;
        RECT  3.070 2.310 3.620 2.730 ;
        RECT  2.900 1.845 3.070 2.730 ;
        RECT  2.350 2.310 2.900 2.730 ;
        RECT  2.180 1.845 2.350 2.730 ;
        RECT  1.785 2.310 2.180 2.730 ;
        RECT  1.615 1.915 1.785 2.730 ;
        RECT  1.095 2.310 1.615 2.730 ;
        RECT  0.835 1.840 1.095 2.730 ;
        RECT  0.330 2.310 0.835 2.730 ;
        RECT  0.160 1.620 0.330 2.730 ;
        RECT  0.000 2.310 0.160 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  2.365 1.050 2.980 1.170 ;
        RECT  2.245 1.050 2.365 1.685 ;
        RECT  1.915 1.050 2.245 1.170 ;
        RECT  1.425 1.565 2.245 1.685 ;
        RECT  1.795 0.625 1.915 1.170 ;
        RECT  0.330 0.625 1.795 0.745 ;
        RECT  1.255 1.565 1.425 1.995 ;
        RECT  0.690 1.565 1.255 1.685 ;
        RECT  0.520 1.565 0.690 1.995 ;
        RECT  0.160 0.535 0.330 0.745 ;
    END
END AND2X8AD
MACRO AND2XLAD
    CLASS CORE ;
    FOREIGN AND2XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.665 1.330 1.805 ;
        END
        AntennaDiffArea 0.149 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.020 0.770 1.375 ;
        END
        AntennaGateArea 0.0424 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.055 0.365 1.315 ;
        RECT  0.070 1.055 0.210 1.655 ;
        END
        AntennaGateArea 0.0424 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.920 -0.210 1.400 0.210 ;
        RECT  0.750 -0.210 0.920 0.660 ;
        RECT  0.000 -0.210 0.750 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.925 2.310 1.400 2.730 ;
        RECT  0.755 1.925 0.925 2.730 ;
        RECT  0.255 2.310 0.755 2.730 ;
        RECT  0.085 1.925 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.920 0.780 1.040 1.615 ;
        RECT  0.270 0.780 0.920 0.900 ;
        RECT  0.390 1.495 0.920 1.615 ;
        RECT  0.100 0.730 0.270 0.900 ;
    END
END AND2XLAD
MACRO AND3X1AD
    CLASS CORE ;
    FOREIGN AND3X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.625 1.610 1.990 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 1.020 1.090 1.375 ;
        END
        AntennaGateArea 0.0474 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 1.020 0.770 1.375 ;
        END
        AntennaGateArea 0.0474 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.145 0.385 1.375 ;
        END
        AntennaGateArea 0.0464 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.205 -0.210 1.680 0.210 ;
        RECT  1.035 -0.210 1.205 0.660 ;
        RECT  0.000 -0.210 1.035 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.195 2.310 1.680 2.730 ;
        RECT  1.025 1.915 1.195 2.730 ;
        RECT  0.615 2.310 1.025 2.730 ;
        RECT  0.445 1.915 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.210 0.780 1.330 1.615 ;
        RECT  0.265 0.780 1.210 0.900 ;
        RECT  0.240 1.495 1.210 1.615 ;
        RECT  0.095 0.710 0.265 0.900 ;
        RECT  0.120 1.495 0.240 2.115 ;
    END
END AND3X1AD
MACRO AND3X2AD
    CLASS CORE ;
    FOREIGN AND3X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.430 1.610 1.990 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 1.020 1.090 1.375 ;
        END
        AntennaGateArea 0.0834 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 1.020 0.770 1.375 ;
        END
        AntennaGateArea 0.0834 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 1.020 0.360 1.375 ;
        RECT  0.070 1.145 0.240 1.375 ;
        END
        AntennaGateArea 0.0834 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.250 -0.210 1.680 0.210 ;
        RECT  0.990 -0.210 1.250 0.650 ;
        RECT  0.000 -0.210 0.990 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.195 2.310 1.680 2.730 ;
        RECT  1.025 2.105 1.195 2.730 ;
        RECT  0.615 2.310 1.025 2.730 ;
        RECT  0.445 1.985 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.210 0.780 1.330 1.615 ;
        RECT  0.265 0.780 1.210 0.900 ;
        RECT  0.265 1.495 1.210 1.615 ;
        RECT  0.095 0.710 0.265 0.900 ;
        RECT  0.145 1.495 0.265 2.155 ;
        RECT  0.095 1.985 0.145 2.155 ;
    END
END AND3X2AD
MACRO AND3X4AD
    CLASS CORE ;
    FOREIGN AND3X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.610 0.725 2.800 1.470 ;
        RECT  2.590 0.725 2.610 2.035 ;
        RECT  2.585 0.725 2.590 0.910 ;
        RECT  2.435 1.315 2.590 2.035 ;
        RECT  2.375 0.375 2.585 0.910 ;
        END
        AntennaDiffArea 0.45 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.270 1.990 1.665 ;
        RECT  0.510 1.545 1.870 1.665 ;
        RECT  0.505 1.145 0.510 1.665 ;
        RECT  0.390 1.040 0.505 1.665 ;
        RECT  0.315 1.040 0.390 1.375 ;
        RECT  0.070 1.145 0.315 1.375 ;
        END
        AntennaGateArea 0.1661 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 1.305 1.750 1.425 ;
        RECT  0.630 0.860 0.810 1.425 ;
        END
        AntennaGateArea 0.1661 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.910 1.375 1.160 ;
        END
        AntennaGateArea 0.1654 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.975 -0.210 3.080 0.210 ;
        RECT  2.785 -0.210 2.975 0.540 ;
        RECT  2.210 -0.210 2.785 0.210 ;
        RECT  2.030 -0.210 2.210 0.675 ;
        RECT  0.380 -0.210 2.030 0.210 ;
        RECT  0.210 -0.210 0.380 0.810 ;
        RECT  0.000 -0.210 0.210 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.950 2.310 3.080 2.730 ;
        RECT  2.785 1.680 2.950 2.730 ;
        RECT  2.175 2.310 2.785 2.730 ;
        RECT  1.305 2.080 2.175 2.730 ;
        RECT  0.715 2.310 1.305 2.730 ;
        RECT  0.455 2.025 0.715 2.730 ;
        RECT  0.000 2.310 0.455 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  2.315 1.030 2.470 1.180 ;
        RECT  2.195 1.030 2.315 1.905 ;
        RECT  1.910 1.030 2.195 1.150 ;
        RECT  0.260 1.785 2.195 1.905 ;
        RECT  1.790 0.620 1.910 1.150 ;
        RECT  1.080 0.620 1.790 0.740 ;
        RECT  0.140 1.510 0.260 2.030 ;
    END
END AND3X4AD
MACRO AND3X6AD
    CLASS CORE ;
    FOREIGN AND3X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.325 0.475 3.495 1.815 ;
        RECT  3.150 0.845 3.325 1.655 ;
        RECT  2.775 1.090 3.150 1.375 ;
        RECT  2.605 0.475 2.775 2.045 ;
        END
        AntennaDiffArea 0.795 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.020 2.120 1.560 ;
        RECT  0.510 1.440 2.000 1.560 ;
        RECT  0.375 1.070 0.510 1.560 ;
        RECT  0.210 1.070 0.375 1.190 ;
        RECT  0.070 0.865 0.210 1.190 ;
        END
        AntennaGateArea 0.2482 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.090 1.840 1.210 ;
        RECT  1.570 0.670 1.690 1.210 ;
        RECT  0.825 0.670 1.570 0.790 ;
        RECT  0.630 0.670 0.825 1.275 ;
        END
        AntennaGateArea 0.2488 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 0.910 1.375 1.170 ;
        END
        AntennaGateArea 0.2488 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.135 -0.210 3.640 0.210 ;
        RECT  2.965 -0.210 3.135 0.675 ;
        RECT  2.345 -0.210 2.965 0.210 ;
        RECT  2.175 -0.210 2.345 0.615 ;
        RECT  0.385 -0.210 2.175 0.210 ;
        RECT  0.190 -0.210 0.385 0.685 ;
        RECT  0.000 -0.210 0.190 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.145 2.310 3.640 2.730 ;
        RECT  2.955 1.865 3.145 2.730 ;
        RECT  2.460 2.310 2.955 2.730 ;
        RECT  2.200 2.010 2.460 2.730 ;
        RECT  1.575 2.310 2.200 2.730 ;
        RECT  0.885 2.165 1.575 2.730 ;
        RECT  0.255 2.310 0.885 2.730 ;
        RECT  0.085 1.475 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  2.405 0.980 2.465 1.240 ;
        RECT  2.285 0.780 2.405 1.800 ;
        RECT  2.010 0.780 2.285 0.900 ;
        RECT  0.400 1.680 2.285 1.800 ;
        RECT  1.890 0.390 2.010 0.900 ;
        RECT  1.100 0.390 1.890 0.510 ;
    END
END AND3X6AD
MACRO AND3X8AD
    CLASS CORE ;
    FOREIGN AND3X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.515 0.620 4.595 1.630 ;
        RECT  4.315 0.475 4.515 2.045 ;
        RECT  4.085 0.620 4.315 1.630 ;
        RECT  3.795 0.620 4.085 0.870 ;
        RECT  3.810 1.380 4.085 1.630 ;
        RECT  3.580 1.380 3.810 2.045 ;
        RECT  3.595 0.440 3.795 0.870 ;
        END
        AntennaDiffArea 0.844 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.050 1.290 3.170 1.620 ;
        RECT  1.550 1.290 3.050 1.410 ;
        RECT  1.190 1.110 1.550 1.410 ;
        RECT  1.030 1.110 1.190 1.230 ;
        END
        AntennaGateArea 0.3326 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.815 1.040 2.985 1.160 ;
        RECT  1.695 0.865 1.815 1.160 ;
        RECT  0.820 0.865 1.695 0.990 ;
        RECT  0.630 0.865 0.820 1.270 ;
        END
        AntennaGateArea 0.3326 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.530 2.770 1.650 ;
        RECT  0.390 1.015 0.510 1.650 ;
        RECT  0.260 1.015 0.390 1.190 ;
        RECT  0.110 0.865 0.260 1.190 ;
        RECT  0.070 0.865 0.110 1.095 ;
        END
        AntennaGateArea 0.3304 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.855 -0.210 5.040 0.210 ;
        RECT  4.735 -0.210 4.855 0.840 ;
        RECT  4.140 -0.210 4.735 0.210 ;
        RECT  3.970 -0.210 4.140 0.415 ;
        RECT  3.455 -0.210 3.970 0.210 ;
        RECT  3.195 -0.210 3.455 0.630 ;
        RECT  1.430 -0.210 3.195 0.210 ;
        RECT  1.170 -0.210 1.430 0.390 ;
        RECT  0.000 -0.210 1.170 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.860 2.310 5.040 2.730 ;
        RECT  4.690 1.845 4.860 2.730 ;
        RECT  4.140 2.310 4.690 2.730 ;
        RECT  3.970 1.845 4.140 2.730 ;
        RECT  3.405 2.310 3.970 2.730 ;
        RECT  2.365 2.130 3.405 2.730 ;
        RECT  1.820 2.310 2.365 2.730 ;
        RECT  1.560 2.020 1.820 2.730 ;
        RECT  1.060 2.310 1.560 2.730 ;
        RECT  0.800 2.020 1.060 2.730 ;
        RECT  0.250 2.310 0.800 2.730 ;
        RECT  0.100 1.480 0.250 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.040 2.520 ;
        LAYER M1 ;
        RECT  3.410 1.000 3.865 1.260 ;
        RECT  3.290 0.750 3.410 1.900 ;
        RECT  3.005 0.750 3.290 0.870 ;
        RECT  0.420 1.780 3.290 1.900 ;
        RECT  2.855 0.515 3.005 0.870 ;
        RECT  2.405 0.515 2.855 0.635 ;
        RECT  2.235 0.385 2.405 0.815 ;
        RECT  0.130 0.515 2.235 0.635 ;
    END
END AND3X8AD
MACRO AND3XLAD
    CLASS CORE ;
    FOREIGN AND3XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.685 1.610 1.805 ;
        END
        AntennaDiffArea 0.143 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 1.020 1.090 1.375 ;
        END
        AntennaGateArea 0.0424 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.555 1.020 0.770 1.375 ;
        END
        AntennaGateArea 0.0424 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.145 0.385 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.205 -0.210 1.680 0.210 ;
        RECT  1.035 -0.210 1.205 0.660 ;
        RECT  0.000 -0.210 1.035 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.195 2.310 1.680 2.730 ;
        RECT  1.025 1.915 1.195 2.730 ;
        RECT  0.615 2.310 1.025 2.730 ;
        RECT  0.445 1.915 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.210 0.780 1.330 1.615 ;
        RECT  0.265 0.780 1.210 0.900 ;
        RECT  0.240 1.495 1.210 1.615 ;
        RECT  0.095 0.730 0.265 0.900 ;
        RECT  0.120 1.495 0.240 2.115 ;
    END
END AND3XLAD
MACRO AND4X1AD
    CLASS CORE ;
    FOREIGN AND4X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.585 2.170 1.960 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.100 0.975 1.600 1.135 ;
        RECT  0.865 0.910 1.100 1.135 ;
        END
        AntennaGateArea 0.0514 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.145 1.905 1.375 2.170 ;
        RECT  0.920 1.905 1.145 2.025 ;
        END
        AntennaGateArea 0.0521 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.770 0.770 1.890 ;
        RECT  0.105 1.740 0.670 1.890 ;
        END
        AntennaGateArea 0.0521 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.990 0.375 1.215 ;
        RECT  0.070 0.990 0.210 1.375 ;
        END
        AntennaGateArea 0.0514 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.800 -0.210 2.240 0.210 ;
        RECT  1.540 -0.210 1.800 0.530 ;
        RECT  0.000 -0.210 1.540 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.755 2.310 2.240 2.730 ;
        RECT  1.585 1.665 1.755 2.730 ;
        RECT  1.040 1.665 1.585 1.785 ;
        RECT  0.255 2.310 1.585 2.730 ;
        RECT  0.920 1.530 1.040 1.785 ;
        RECT  0.775 1.530 0.920 1.650 ;
        RECT  0.085 2.010 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.770 0.650 1.890 1.410 ;
        RECT  0.325 0.650 1.770 0.780 ;
        RECT  1.420 1.290 1.770 1.410 ;
        RECT  1.160 1.290 1.420 1.545 ;
        RECT  0.615 1.290 1.160 1.410 ;
        RECT  0.495 1.290 0.615 1.570 ;
        RECT  0.435 1.400 0.495 1.570 ;
        RECT  0.155 0.650 0.325 0.820 ;
    END
END AND4X1AD
MACRO AND4X2AD
    CLASS CORE ;
    FOREIGN AND4X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.430 2.170 1.960 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.100 1.020 1.600 1.140 ;
        RECT  0.865 0.910 1.100 1.140 ;
        END
        AntennaGateArea 0.0904 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.145 1.905 1.375 2.170 ;
        RECT  0.920 1.905 1.145 2.025 ;
        END
        AntennaGateArea 0.09 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.740 0.770 1.980 ;
        RECT  0.105 1.740 0.510 1.890 ;
        END
        AntennaGateArea 0.09 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.045 0.375 1.215 ;
        RECT  0.070 1.045 0.210 1.375 ;
        END
        AntennaGateArea 0.0904 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.210 2.240 0.210 ;
        RECT  1.555 -0.210 1.725 0.530 ;
        RECT  0.000 -0.210 1.555 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.755 2.310 2.240 2.730 ;
        RECT  1.585 1.665 1.755 2.730 ;
        RECT  1.040 1.665 1.585 1.785 ;
        RECT  0.255 2.310 1.585 2.730 ;
        RECT  0.920 1.500 1.040 1.785 ;
        RECT  0.775 1.500 0.920 1.620 ;
        RECT  0.085 2.010 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.770 0.650 1.890 1.380 ;
        RECT  0.325 0.650 1.770 0.780 ;
        RECT  1.420 1.260 1.770 1.380 ;
        RECT  1.160 1.260 1.420 1.545 ;
        RECT  0.615 1.260 1.160 1.380 ;
        RECT  0.495 1.260 0.615 1.570 ;
        RECT  0.435 1.400 0.495 1.570 ;
        RECT  0.155 0.475 0.325 0.905 ;
    END
END AND4X2AD
MACRO AND4X4AD
    CLASS CORE ;
    FOREIGN AND4X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.200 0.715 3.290 1.565 ;
        RECT  3.155 0.415 3.200 1.565 ;
        RECT  3.150 0.415 3.155 1.865 ;
        RECT  3.025 0.415 3.150 0.845 ;
        RECT  2.985 1.435 3.150 1.865 ;
        END
        AntennaDiffArea 0.45 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.385 1.020 2.505 1.730 ;
        RECT  0.210 1.610 2.385 1.730 ;
        RECT  0.070 1.425 0.210 1.935 ;
        END
        AntennaGateArea 0.1795 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.085 1.200 2.205 1.490 ;
        RECT  0.490 1.370 2.085 1.490 ;
        RECT  0.350 0.865 0.490 1.490 ;
        END
        AntennaGateArea 0.179 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 0.670 1.895 1.250 ;
        RECT  0.770 0.670 1.775 0.790 ;
        RECT  0.770 1.070 1.010 1.190 ;
        RECT  0.630 0.670 0.770 1.190 ;
        END
        AntennaGateArea 0.179 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.145 0.910 1.655 1.150 ;
        END
        AntennaGateArea 0.179 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.555 -0.210 3.640 0.210 ;
        RECT  3.385 -0.210 3.555 0.595 ;
        RECT  2.725 -0.210 3.385 0.210 ;
        RECT  2.555 -0.210 2.725 0.615 ;
        RECT  0.230 -0.210 2.555 0.210 ;
        RECT  0.110 -0.210 0.230 0.880 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.515 2.310 3.640 2.730 ;
        RECT  3.345 1.730 3.515 2.730 ;
        RECT  2.725 2.310 3.345 2.730 ;
        RECT  2.555 2.105 2.725 2.730 ;
        RECT  1.960 2.310 2.555 2.730 ;
        RECT  1.790 2.105 1.960 2.730 ;
        RECT  1.265 2.310 1.790 2.730 ;
        RECT  1.005 1.870 1.265 2.730 ;
        RECT  0.000 2.310 1.005 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  2.805 1.010 3.005 1.270 ;
        RECT  2.685 0.780 2.805 1.970 ;
        RECT  2.225 0.780 2.685 0.900 ;
        RECT  1.385 1.850 2.685 1.970 ;
        RECT  2.105 0.430 2.225 0.900 ;
        RECT  1.200 0.430 2.105 0.550 ;
    END
END AND4X4AD
MACRO AND4X6AD
    CLASS CORE ;
    FOREIGN AND4X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.775 0.475 4.945 0.910 ;
        RECT  4.775 1.475 4.945 1.935 ;
        RECT  4.730 0.730 4.775 0.910 ;
        RECT  4.730 1.475 4.775 1.655 ;
        RECT  4.550 0.730 4.730 1.655 ;
        RECT  4.225 0.730 4.550 0.910 ;
        RECT  4.225 1.475 4.550 1.655 ;
        RECT  4.055 0.415 4.225 0.910 ;
        RECT  4.055 1.475 4.225 1.970 ;
        END
        AntennaDiffArea 0.795 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.570 0.990 3.690 1.880 ;
        RECT  1.350 1.760 3.570 1.880 ;
        RECT  1.190 1.145 1.350 1.880 ;
        END
        AntennaGateArea 0.2688 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.320 1.320 3.440 1.640 ;
        RECT  1.890 1.520 3.320 1.640 ;
        RECT  1.745 0.865 1.890 1.640 ;
        RECT  1.050 0.865 1.745 0.985 ;
        RECT  0.930 0.865 1.050 1.260 ;
        END
        AntennaGateArea 0.269 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.250 1.280 3.160 1.400 ;
        RECT  2.130 0.625 2.250 1.400 ;
        RECT  0.770 0.625 2.130 0.745 ;
        RECT  0.620 0.625 0.770 1.375 ;
        END
        AntennaGateArea 0.2684 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 1.030 2.650 1.150 ;
        RECT  2.370 0.385 2.490 1.150 ;
        RECT  0.490 0.385 2.370 0.505 ;
        RECT  0.370 0.385 0.490 1.375 ;
        RECT  0.320 0.865 0.370 1.375 ;
        END
        AntennaGateArea 0.2688 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.630 -0.210 5.040 0.210 ;
        RECT  4.370 -0.210 4.630 0.560 ;
        RECT  3.910 -0.210 4.370 0.210 ;
        RECT  3.650 -0.210 3.910 0.560 ;
        RECT  1.590 -0.210 3.650 0.210 ;
        RECT  1.330 -0.210 1.590 0.265 ;
        RECT  0.000 -0.210 1.330 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.585 2.310 5.040 2.730 ;
        RECT  4.415 1.905 4.585 2.730 ;
        RECT  3.795 2.310 4.415 2.730 ;
        RECT  3.625 2.245 3.795 2.730 ;
        RECT  2.880 2.310 3.625 2.730 ;
        RECT  2.710 2.245 2.880 2.730 ;
        RECT  2.120 2.310 2.710 2.730 ;
        RECT  1.950 2.245 2.120 2.730 ;
        RECT  1.360 2.310 1.950 2.730 ;
        RECT  1.190 2.245 1.360 2.730 ;
        RECT  0.615 2.310 1.190 2.730 ;
        RECT  0.445 1.850 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.040 2.520 ;
        LAYER M1 ;
        RECT  3.930 1.085 4.410 1.205 ;
        RECT  3.810 0.680 3.930 2.125 ;
        RECT  2.730 0.680 3.810 0.800 ;
        RECT  0.980 2.005 3.810 2.125 ;
        RECT  2.610 0.485 2.730 0.800 ;
        RECT  0.835 1.560 0.980 2.125 ;
        RECT  0.810 1.560 0.835 2.105 ;
        RECT  0.190 1.560 0.810 1.680 ;
        RECT  0.190 0.450 0.230 0.710 ;
        RECT  0.070 0.450 0.190 1.680 ;
    END
END AND4X6AD
MACRO AND4X8AD
    CLASS CORE ;
    FOREIGN AND4X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.760 0.430 6.020 1.980 ;
        RECT  5.530 0.665 5.760 1.600 ;
        RECT  5.325 0.665 5.530 0.915 ;
        RECT  5.280 1.350 5.530 1.600 ;
        RECT  5.110 0.370 5.325 0.915 ;
        RECT  5.110 1.350 5.280 2.045 ;
        END
        AntennaDiffArea 0.844 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.630 0.980 4.750 1.860 ;
        RECT  2.450 1.740 4.630 1.860 ;
        RECT  2.310 1.190 2.450 1.860 ;
        RECT  0.350 1.740 2.310 1.860 ;
        END
        AntennaGateArea 0.3606 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.310 1.200 4.430 1.620 ;
        RECT  2.920 1.500 4.310 1.620 ;
        RECT  2.800 1.145 2.920 1.620 ;
        RECT  2.710 1.145 2.800 1.375 ;
        RECT  2.590 0.900 2.710 1.375 ;
        RECT  2.070 0.900 2.590 1.020 ;
        RECT  1.950 0.900 2.070 1.620 ;
        RECT  0.630 1.500 1.950 1.620 ;
        RECT  0.510 1.330 0.630 1.620 ;
        END
        AntennaGateArea 0.3601 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.270 1.260 4.060 1.380 ;
        RECT  3.090 0.905 3.270 1.380 ;
        RECT  2.950 0.905 3.090 1.025 ;
        RECT  2.830 0.660 2.950 1.025 ;
        RECT  1.820 0.660 2.830 0.780 ;
        RECT  1.700 0.660 1.820 1.375 ;
        RECT  1.470 1.145 1.700 1.375 ;
        END
        AntennaGateArea 0.3606 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.665 3.570 1.140 ;
        RECT  3.190 0.665 3.450 0.785 ;
        RECT  3.070 0.420 3.190 0.785 ;
        RECT  1.580 0.420 3.070 0.540 ;
        RECT  1.460 0.420 1.580 0.985 ;
        RECT  1.330 0.865 1.460 0.985 ;
        RECT  1.030 0.865 1.330 1.095 ;
        END
        AntennaGateArea 0.3606 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.335 -0.210 6.440 0.210 ;
        RECT  6.165 -0.210 6.335 0.785 ;
        RECT  5.615 -0.210 6.165 0.210 ;
        RECT  5.445 -0.210 5.615 0.525 ;
        RECT  4.940 -0.210 5.445 0.210 ;
        RECT  4.680 -0.210 4.940 0.510 ;
        RECT  2.610 -0.210 4.680 0.210 ;
        RECT  2.350 -0.210 2.610 0.300 ;
        RECT  0.230 -0.210 2.350 0.210 ;
        RECT  0.110 -0.210 0.230 0.790 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.335 2.310 6.440 2.730 ;
        RECT  6.165 1.735 6.335 2.730 ;
        RECT  5.615 2.310 6.165 2.730 ;
        RECT  5.445 1.735 5.615 2.730 ;
        RECT  4.770 2.310 5.445 2.730 ;
        RECT  4.600 2.220 4.770 2.730 ;
        RECT  3.875 2.310 4.600 2.730 ;
        RECT  3.705 2.220 3.875 2.730 ;
        RECT  3.115 2.310 3.705 2.730 ;
        RECT  2.945 2.220 3.115 2.730 ;
        RECT  2.355 2.310 2.945 2.730 ;
        RECT  2.185 2.220 2.355 2.730 ;
        RECT  1.595 2.310 2.185 2.730 ;
        RECT  1.425 2.220 1.595 2.730 ;
        RECT  0.000 2.310 1.425 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.440 2.520 ;
        LAYER M1 ;
        RECT  4.990 1.085 5.410 1.205 ;
        RECT  4.870 0.670 4.990 2.100 ;
        RECT  4.000 0.670 4.870 0.790 ;
        RECT  0.230 1.980 4.870 2.100 ;
        RECT  3.880 0.425 4.000 0.790 ;
        RECT  3.530 0.425 3.880 0.545 ;
        RECT  1.220 0.470 1.340 0.730 ;
        RECT  0.640 0.610 1.220 0.730 ;
        RECT  0.520 0.610 0.640 1.210 ;
        RECT  0.230 1.090 0.520 1.210 ;
        RECT  0.110 1.090 0.230 2.100 ;
    END
END AND4X8AD
MACRO AND4XLAD
    CLASS CORE ;
    FOREIGN AND4XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.585 2.170 1.730 ;
        END
        AntennaDiffArea 0.155 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.100 0.975 1.600 1.135 ;
        RECT  0.865 0.910 1.100 1.135 ;
        END
        AntennaGateArea 0.0424 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.145 1.905 1.375 2.170 ;
        RECT  0.920 1.905 1.145 2.025 ;
        END
        AntennaGateArea 0.0431 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.770 0.770 1.890 ;
        RECT  0.105 1.740 0.670 1.890 ;
        END
        AntennaGateArea 0.0431 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.990 0.375 1.215 ;
        RECT  0.070 0.990 0.210 1.375 ;
        END
        AntennaGateArea 0.0424 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.800 -0.210 2.240 0.210 ;
        RECT  1.540 -0.210 1.800 0.530 ;
        RECT  0.000 -0.210 1.540 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.755 2.310 2.240 2.730 ;
        RECT  1.585 1.590 1.755 2.730 ;
        RECT  1.040 1.665 1.585 1.785 ;
        RECT  0.255 2.310 1.585 2.730 ;
        RECT  0.920 1.530 1.040 1.785 ;
        RECT  0.775 1.530 0.920 1.650 ;
        RECT  0.085 2.010 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.770 0.650 1.890 1.410 ;
        RECT  0.325 0.650 1.770 0.780 ;
        RECT  1.420 1.290 1.770 1.410 ;
        RECT  1.160 1.290 1.420 1.545 ;
        RECT  0.615 1.290 1.160 1.410 ;
        RECT  0.495 1.290 0.615 1.570 ;
        RECT  0.435 1.400 0.495 1.570 ;
        RECT  0.155 0.650 0.325 0.820 ;
    END
END AND4XLAD
MACRO ANTENNAAD
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNAAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.535 0.585 0.625 0.815 ;
        RECT  0.305 0.585 0.535 1.965 ;
        RECT  0.070 0.585 0.305 0.815 ;
        END
        AntennaDiffArea 0.663 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.210 0.840 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.310 0.840 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 0.840 2.520 ;
	 END
END ANTENNAAD
MACRO AO21X1AD
    CLASS CORE ;
    FOREIGN AO21X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.865 0.520 1.890 1.595 ;
        RECT  1.750 0.520 1.865 1.920 ;
        RECT  1.530 0.520 1.750 0.640 ;
        RECT  1.695 1.490 1.750 1.920 ;
        END
        AntennaDiffArea 0.221 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.895 1.030 1.145 1.375 ;
        END
        AntennaGateArea 0.0464 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.975 0.370 1.235 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.0464 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.540 1.030 0.770 1.375 ;
        END
        AntennaGateArea 0.0464 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.370 -0.210 1.960 0.210 ;
        RECT  1.110 -0.210 1.370 0.670 ;
        RECT  0.265 -0.210 1.110 0.210 ;
        RECT  0.095 -0.210 0.265 0.745 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.505 2.310 1.960 2.730 ;
        RECT  1.335 1.830 1.505 2.730 ;
        RECT  0.590 2.310 1.335 2.730 ;
        RECT  0.330 1.495 0.590 2.730 ;
        RECT  0.000 2.310 0.330 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.450 0.980 1.570 1.240 ;
        RECT  1.330 0.790 1.450 1.615 ;
        RECT  0.885 0.790 1.330 0.910 ;
        RECT  1.000 1.495 1.330 1.615 ;
        RECT  0.715 0.575 0.885 0.910 ;
    END
END AO21X1AD
MACRO AO21X2AD
    CLASS CORE ;
    FOREIGN AO21X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.875 0.710 1.890 1.680 ;
        RECT  1.750 0.710 1.875 1.990 ;
        RECT  1.720 0.710 1.750 0.850 ;
        RECT  1.705 1.560 1.750 1.990 ;
        RECT  1.600 0.330 1.720 0.850 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.895 1.020 1.125 1.375 ;
        END
        AntennaGateArea 0.0744 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 1.010 0.395 1.375 ;
        RECT  0.070 1.145 0.190 1.375 ;
        END
        AntennaGateArea 0.0844 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.540 1.020 0.770 1.375 ;
        END
        AntennaGateArea 0.0844 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.430 -0.210 1.960 0.210 ;
        RECT  1.170 -0.210 1.430 0.650 ;
        RECT  0.265 -0.210 1.170 0.210 ;
        RECT  0.095 -0.210 0.265 0.875 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 2.310 1.960 2.730 ;
        RECT  1.345 1.945 1.515 2.730 ;
        RECT  0.545 2.310 1.345 2.730 ;
        RECT  0.375 1.510 0.545 2.730 ;
        RECT  0.000 2.310 0.375 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.450 1.000 1.605 1.260 ;
        RECT  1.330 0.770 1.450 1.615 ;
        RECT  0.885 0.770 1.330 0.890 ;
        RECT  1.000 1.495 1.330 1.615 ;
        RECT  0.715 0.680 0.885 0.890 ;
    END
END AO21X2AD
MACRO AO21X4AD
    CLASS CORE ;
    FOREIGN AO21X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.795 2.450 1.515 ;
        RECT  2.075 0.795 2.310 0.935 ;
        RECT  2.075 1.375 2.310 1.515 ;
        RECT  1.905 0.375 2.075 0.935 ;
        RECT  1.905 1.375 2.075 1.995 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 1.000 1.090 1.375 ;
        END
        AntennaGateArea 0.147 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.005 0.420 1.265 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 1.000 0.770 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 -0.210 2.520 0.210 ;
        RECT  2.265 -0.210 2.435 0.675 ;
        RECT  1.440 -0.210 2.265 0.210 ;
        RECT  1.440 0.445 1.640 0.565 ;
        RECT  1.320 -0.210 1.440 0.565 ;
        RECT  0.270 -0.210 1.320 0.210 ;
        RECT  1.120 0.445 1.320 0.565 ;
        RECT  0.100 -0.210 0.270 0.735 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 2.310 2.520 2.730 ;
        RECT  2.265 1.725 2.435 2.730 ;
        RECT  1.715 2.310 2.265 2.730 ;
        RECT  1.545 1.570 1.715 2.730 ;
        RECT  0.645 2.310 1.545 2.730 ;
        RECT  0.475 1.845 0.645 2.730 ;
        RECT  0.000 2.310 0.475 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.375 1.065 2.180 1.235 ;
        RECT  1.255 0.750 1.375 1.995 ;
        RECT  0.895 0.750 1.255 0.870 ;
        RECT  1.205 1.565 1.255 1.995 ;
        RECT  0.845 1.495 1.015 1.995 ;
        RECT  0.725 0.395 0.895 0.870 ;
        RECT  0.270 1.495 0.845 1.615 ;
        RECT  0.100 1.495 0.270 1.995 ;
    END
END AO21X4AD
MACRO AO21XLAD
    CLASS CORE ;
    FOREIGN AO21XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.715 1.890 1.915 ;
        RECT  1.575 0.715 1.750 0.885 ;
        RECT  1.705 1.745 1.750 1.915 ;
        END
        AntennaDiffArea 0.148 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.895 1.030 1.125 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 1.010 0.395 1.375 ;
        RECT  0.070 1.145 0.190 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.530 1.030 0.770 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.370 -0.210 1.960 0.210 ;
        RECT  1.110 -0.210 1.370 0.670 ;
        RECT  0.265 -0.210 1.110 0.210 ;
        RECT  0.095 -0.210 0.265 0.885 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.505 2.310 1.960 2.730 ;
        RECT  1.335 1.845 1.505 2.730 ;
        RECT  0.590 2.310 1.335 2.730 ;
        RECT  0.330 1.495 0.590 2.730 ;
        RECT  0.000 2.310 0.330 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.450 1.005 1.625 1.455 ;
        RECT  1.330 0.790 1.450 1.615 ;
        RECT  0.885 0.790 1.330 0.910 ;
        RECT  1.020 1.495 1.330 1.615 ;
        RECT  0.715 0.715 0.885 0.910 ;
    END
END AO21XLAD
MACRO AO22X1AD
    CLASS CORE ;
    FOREIGN AO22X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.155 0.505 2.170 1.655 ;
        RECT  2.030 0.505 2.155 1.955 ;
        RECT  1.855 0.505 2.030 0.765 ;
        RECT  1.985 1.525 2.030 1.955 ;
        END
        AntennaDiffArea 0.218 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.990 0.370 1.250 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.540 0.860 0.770 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.865 1.385 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 0.865 1.070 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.610 -0.210 2.240 0.210 ;
        RECT  1.350 -0.210 1.610 0.465 ;
        RECT  0.265 -0.210 1.350 0.210 ;
        RECT  0.095 -0.210 0.265 0.745 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.820 2.310 2.240 2.730 ;
        RECT  1.560 2.220 1.820 2.730 ;
        RECT  0.590 2.310 1.560 2.730 ;
        RECT  0.330 1.500 0.590 2.730 ;
        RECT  0.000 2.310 0.330 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.615 0.600 1.735 1.620 ;
        RECT  0.660 0.600 1.615 0.720 ;
        RECT  1.000 1.500 1.615 1.620 ;
    END
END AO22X1AD
MACRO AO22X2AD
    CLASS CORE ;
    FOREIGN AO22X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.410 1.140 2.450 1.375 ;
        RECT  2.270 0.355 2.410 2.030 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.985 0.380 1.245 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.083 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 0.855 0.770 1.375 ;
        END
        AntennaGateArea 0.0835 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 0.855 1.610 1.375 ;
        END
        AntennaGateArea 0.0835 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.855 1.100 1.375 ;
        END
        AntennaGateArea 0.0835 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.840 -0.210 2.520 0.210 ;
        RECT  1.840 0.375 1.990 0.495 ;
        RECT  1.640 -0.210 1.840 0.495 ;
        RECT  0.255 -0.210 1.640 0.210 ;
        RECT  1.470 0.375 1.640 0.495 ;
        RECT  0.085 -0.210 0.255 0.675 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.075 2.310 2.520 2.730 ;
        RECT  1.905 1.790 2.075 2.730 ;
        RECT  0.660 2.310 1.905 2.730 ;
        RECT  0.400 1.735 0.660 2.730 ;
        RECT  0.000 2.310 0.400 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.030 0.615 2.150 1.615 ;
        RECT  0.905 0.615 2.030 0.735 ;
        RECT  1.120 1.495 2.030 1.615 ;
        RECT  0.975 1.735 1.740 1.855 ;
        RECT  0.805 1.495 0.975 1.855 ;
        RECT  0.735 0.480 0.905 0.735 ;
        RECT  0.255 1.495 0.805 1.615 ;
        RECT  0.085 1.495 0.255 1.765 ;
    END
END AO22X2AD
MACRO AO22X4AD
    CLASS CORE ;
    FOREIGN AO22X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.775 2.730 1.535 ;
        RECT  2.355 0.775 2.590 0.905 ;
        RECT  2.355 1.405 2.590 1.535 ;
        RECT  2.185 0.355 2.355 0.905 ;
        RECT  2.185 1.405 2.355 1.980 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 1.010 0.475 1.375 ;
        RECT  0.070 1.145 0.305 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 0.995 0.790 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 0.995 1.610 1.375 ;
        END
        AntennaGateArea 0.1629 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.995 1.200 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.715 -0.210 2.800 0.210 ;
        RECT  2.545 -0.210 2.715 0.635 ;
        RECT  1.845 -0.210 2.545 0.210 ;
        RECT  1.845 0.490 2.010 0.610 ;
        RECT  1.675 -0.210 1.845 0.610 ;
        RECT  0.350 -0.210 1.675 0.210 ;
        RECT  1.490 0.490 1.675 0.610 ;
        RECT  0.180 -0.210 0.350 0.810 ;
        RECT  0.000 -0.210 0.180 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.715 2.310 2.800 2.730 ;
        RECT  2.545 1.655 2.715 2.730 ;
        RECT  1.995 2.310 2.545 2.730 ;
        RECT  1.825 2.105 1.995 2.730 ;
        RECT  0.615 2.310 1.825 2.730 ;
        RECT  0.445 1.735 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  1.910 1.025 2.450 1.285 ;
        RECT  1.790 0.755 1.910 1.615 ;
        RECT  1.005 0.755 1.790 0.875 ;
        RECT  1.335 1.495 1.790 1.615 ;
        RECT  1.525 1.735 1.695 2.060 ;
        RECT  0.975 1.940 1.525 2.060 ;
        RECT  1.165 1.495 1.335 1.795 ;
        RECT  0.835 0.390 1.005 0.875 ;
        RECT  0.805 1.495 0.975 2.060 ;
        RECT  0.255 1.495 0.805 1.615 ;
        RECT  0.085 1.495 0.255 1.950 ;
    END
END AO22X4AD
MACRO AO22XLAD
    CLASS CORE ;
    FOREIGN AO22XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.575 2.170 1.980 ;
        RECT  1.975 0.575 2.030 0.745 ;
        RECT  1.965 1.810 2.030 1.980 ;
        END
        AntennaDiffArea 0.14 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.865 0.410 1.190 ;
        RECT  0.070 0.865 0.210 1.095 ;
        END
        AntennaGateArea 0.0404 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 0.865 0.770 1.280 ;
        END
        AntennaGateArea 0.0404 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 0.865 1.610 1.260 ;
        END
        AntennaGateArea 0.04 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 0.865 1.070 1.280 ;
        END
        AntennaGateArea 0.04 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.735 -0.210 2.240 0.210 ;
        RECT  1.475 -0.210 1.735 0.505 ;
        RECT  0.285 -0.210 1.475 0.210 ;
        RECT  0.115 -0.210 0.285 0.745 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.775 2.310 2.240 2.730 ;
        RECT  1.605 1.905 1.775 2.730 ;
        RECT  0.665 2.310 1.605 2.730 ;
        RECT  0.495 1.805 0.665 2.730 ;
        RECT  0.000 2.310 0.495 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.855 0.980 1.900 1.240 ;
        RECT  1.735 0.625 1.855 1.240 ;
        RECT  1.645 1.400 1.785 1.520 ;
        RECT  1.310 0.625 1.735 0.745 ;
        RECT  1.525 1.400 1.645 1.785 ;
        RECT  1.020 1.665 1.525 1.785 ;
        RECT  1.310 1.375 1.360 1.545 ;
        RECT  1.190 0.625 1.310 1.545 ;
        RECT  0.925 0.625 1.190 0.745 ;
        RECT  0.900 1.400 1.020 1.785 ;
        RECT  0.755 0.575 0.925 0.745 ;
        RECT  0.070 1.400 0.900 1.520 ;
    END
END AO22XLAD
MACRO AO2B2BX1AD
    CLASS CORE ;
    FOREIGN AO2B2BX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.265 0.630 3.290 1.595 ;
        RECT  3.150 0.630 3.265 1.880 ;
        RECT  3.095 0.630 3.150 0.800 ;
        RECT  3.095 1.450 3.150 1.880 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN B1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 1.025 0.350 1.285 ;
        RECT  0.070 0.865 0.230 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B1N
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.865 1.340 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.865 2.730 1.240 ;
        RECT  2.475 0.980 2.590 1.240 ;
        END
        AntennaGateArea 0.0403 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.460 0.865 1.650 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.930 -0.210 3.360 0.210 ;
        RECT  2.670 -0.210 2.930 0.325 ;
        RECT  2.210 -0.210 2.670 0.210 ;
        RECT  1.950 -0.210 2.210 0.330 ;
        RECT  0.880 -0.210 1.950 0.210 ;
        RECT  0.710 -0.210 0.880 0.770 ;
        RECT  0.000 -0.210 0.710 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.905 2.310 3.360 2.730 ;
        RECT  2.735 1.455 2.905 2.730 ;
        RECT  1.240 2.310 2.735 2.730 ;
        RECT  0.980 1.500 1.240 2.730 ;
        RECT  0.255 2.310 0.980 2.730 ;
        RECT  0.085 1.915 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.970 1.005 3.030 1.265 ;
        RECT  2.850 0.455 2.970 1.265 ;
        RECT  1.910 0.455 2.850 0.575 ;
        RECT  2.150 1.400 2.550 1.520 ;
        RECT  2.150 0.695 2.470 0.815 ;
        RECT  2.030 0.695 2.150 1.520 ;
        RECT  1.790 0.455 1.910 1.620 ;
        RECT  1.275 0.625 1.790 0.745 ;
        RECT  1.650 1.500 1.790 1.620 ;
        RECT  0.590 1.020 1.005 1.280 ;
        RECT  0.470 0.625 0.590 1.620 ;
        RECT  0.125 0.625 0.470 0.745 ;
        RECT  0.330 1.500 0.470 1.620 ;
    END
END AO2B2BX1AD
MACRO AO2B2BX2AD
    CLASS CORE ;
    FOREIGN AO2B2BX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.265 0.665 3.290 1.615 ;
        RECT  3.150 0.370 3.265 2.160 ;
        RECT  3.095 0.370 3.150 0.800 ;
        RECT  3.095 1.470 3.150 2.160 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN B1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 1.020 0.330 1.280 ;
        RECT  0.070 0.865 0.230 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END B1N
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.865 1.340 1.375 ;
        END
        AntennaGateArea 0.0834 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.455 1.065 2.730 1.375 ;
        END
        AntennaGateArea 0.0603 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.865 1.660 1.375 ;
        END
        AntennaGateArea 0.0834 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.950 -0.210 3.360 0.210 ;
        RECT  2.690 -0.210 2.950 0.390 ;
        RECT  2.210 -0.210 2.690 0.210 ;
        RECT  1.950 -0.210 2.210 0.400 ;
        RECT  0.880 -0.210 1.950 0.210 ;
        RECT  0.710 -0.210 0.880 0.840 ;
        RECT  0.000 -0.210 0.710 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.905 2.310 3.360 2.730 ;
        RECT  2.735 1.585 2.905 2.730 ;
        RECT  1.240 2.310 2.735 2.730 ;
        RECT  0.980 1.500 1.240 2.730 ;
        RECT  0.255 2.310 0.980 2.730 ;
        RECT  0.085 2.000 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.970 1.005 3.030 1.265 ;
        RECT  2.850 0.520 2.970 1.265 ;
        RECT  1.900 0.520 2.850 0.640 ;
        RECT  2.140 0.760 2.550 0.880 ;
        RECT  2.140 1.500 2.550 1.620 ;
        RECT  2.020 0.760 2.140 1.620 ;
        RECT  1.780 0.520 1.900 1.680 ;
        RECT  1.275 0.620 1.780 0.740 ;
        RECT  1.695 1.510 1.780 1.680 ;
        RECT  0.590 1.020 1.005 1.280 ;
        RECT  0.470 0.565 0.590 1.615 ;
        RECT  0.170 0.565 0.470 0.735 ;
        RECT  0.330 1.495 0.470 1.615 ;
    END
END AO2B2BX2AD
MACRO AO2B2BX4AD
    CLASS CORE ;
    FOREIGN AO2B2BX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.455 0.390 3.570 1.615 ;
        RECT  3.430 0.390 3.455 2.165 ;
        RECT  3.285 0.390 3.430 0.820 ;
        RECT  3.285 1.475 3.430 2.165 ;
        END
        AntennaDiffArea 0.47 ;
    END Y
    PIN B1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 1.020 0.370 1.280 ;
        RECT  0.120 1.020 0.300 1.375 ;
        RECT  0.070 1.145 0.120 1.375 ;
        END
        AntennaGateArea 0.0674 ;
    END B1N
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.865 1.440 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 1.015 2.830 1.330 ;
        END
        AntennaGateArea 0.0674 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.740 0.865 1.890 1.275 ;
        RECT  1.580 1.000 1.740 1.275 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.810 -0.210 3.920 0.210 ;
        RECT  3.690 -0.210 3.810 0.865 ;
        RECT  3.130 -0.210 3.690 0.210 ;
        RECT  2.870 -0.210 3.130 0.390 ;
        RECT  2.275 -0.210 2.870 0.210 ;
        RECT  2.015 -0.210 2.275 0.390 ;
        RECT  0.840 -0.210 2.015 0.210 ;
        RECT  0.840 0.525 1.015 0.645 ;
        RECT  0.640 -0.210 0.840 0.645 ;
        RECT  0.000 -0.210 0.640 0.210 ;
        RECT  0.495 0.525 0.640 0.645 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.810 2.310 3.920 2.730 ;
        RECT  3.690 1.500 3.810 2.730 ;
        RECT  3.085 2.310 3.690 2.730 ;
        RECT  2.915 1.995 3.085 2.730 ;
        RECT  1.205 2.310 2.915 2.730 ;
        RECT  1.035 1.770 1.205 2.730 ;
        RECT  0.255 2.310 1.035 2.730 ;
        RECT  0.085 2.000 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  3.160 1.005 3.280 1.265 ;
        RECT  3.040 0.520 3.160 1.840 ;
        RECT  1.650 0.520 3.040 0.640 ;
        RECT  1.975 1.720 3.040 1.840 ;
        RECT  2.425 0.760 2.750 0.880 ;
        RECT  2.425 1.450 2.750 1.570 ;
        RECT  2.305 0.760 2.425 1.570 ;
        RECT  1.600 1.970 2.390 2.090 ;
        RECT  2.035 1.020 2.305 1.280 ;
        RECT  1.805 1.410 1.975 1.840 ;
        RECT  1.390 0.340 1.650 0.720 ;
        RECT  1.430 1.495 1.600 2.090 ;
        RECT  0.870 1.495 1.430 1.615 ;
        RECT  0.630 1.065 1.070 1.235 ;
        RECT  0.750 1.495 0.870 2.095 ;
        RECT  0.660 1.925 0.750 2.095 ;
        RECT  0.510 0.780 0.630 1.610 ;
        RECT  0.305 0.780 0.510 0.900 ;
        RECT  0.345 1.490 0.510 1.610 ;
        RECT  0.135 0.695 0.305 0.900 ;
    END
END AO2B2BX4AD
MACRO AO2B2BXLAD
    CLASS CORE ;
    FOREIGN AO2B2BXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.670 3.290 1.675 ;
        RECT  3.095 0.670 3.150 0.840 ;
        RECT  3.095 1.505 3.150 1.675 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN B1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.000 0.370 1.260 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B1N
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.865 1.340 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.865 2.730 1.255 ;
        RECT  2.475 0.995 2.590 1.255 ;
        END
        AntennaGateArea 0.0404 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 0.865 1.630 1.280 ;
        RECT  1.470 0.865 1.610 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.930 -0.210 3.360 0.210 ;
        RECT  2.670 -0.210 2.930 0.330 ;
        RECT  2.180 -0.210 2.670 0.210 ;
        RECT  1.920 -0.210 2.180 0.330 ;
        RECT  0.850 -0.210 1.920 0.210 ;
        RECT  0.730 -0.210 0.850 0.815 ;
        RECT  0.000 -0.210 0.730 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.905 2.310 3.360 2.730 ;
        RECT  2.735 1.480 2.905 2.730 ;
        RECT  1.240 2.310 2.735 2.730 ;
        RECT  0.980 1.500 1.240 2.730 ;
        RECT  0.255 2.310 0.980 2.730 ;
        RECT  0.085 1.915 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.970 0.995 3.030 1.255 ;
        RECT  2.850 0.455 2.970 1.255 ;
        RECT  1.870 0.455 2.850 0.575 ;
        RECT  2.110 1.400 2.550 1.520 ;
        RECT  2.110 0.695 2.470 0.815 ;
        RECT  1.990 0.695 2.110 1.520 ;
        RECT  1.750 0.455 1.870 1.645 ;
        RECT  1.275 0.625 1.750 0.745 ;
        RECT  1.695 1.475 1.750 1.645 ;
        RECT  0.610 1.065 1.000 1.235 ;
        RECT  0.490 0.625 0.610 1.620 ;
        RECT  0.125 0.625 0.490 0.745 ;
        RECT  0.330 1.500 0.490 1.620 ;
    END
END AO2B2BXLAD
MACRO AO2B2X1AD
    CLASS CORE ;
    FOREIGN AO2B2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.705 0.630 2.730 1.540 ;
        RECT  2.590 0.630 2.705 1.880 ;
        RECT  2.535 0.630 2.590 0.800 ;
        RECT  2.535 1.450 2.590 1.880 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 0.960 0.430 1.375 ;
        RECT  0.070 1.145 0.230 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.960 0.770 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.865 2.170 1.245 ;
        RECT  1.915 0.975 2.030 1.245 ;
        END
        AntennaGateArea 0.0403 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 0.960 1.090 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.370 -0.210 2.800 0.210 ;
        RECT  2.110 -0.210 2.370 0.330 ;
        RECT  1.585 -0.210 2.110 0.210 ;
        RECT  1.325 -0.210 1.585 0.330 ;
        RECT  0.270 -0.210 1.325 0.210 ;
        RECT  0.100 -0.210 0.270 0.840 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.345 2.310 2.800 2.730 ;
        RECT  2.175 1.455 2.345 2.730 ;
        RECT  0.610 2.310 2.175 2.730 ;
        RECT  0.350 1.500 0.610 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.410 1.005 2.470 1.265 ;
        RECT  2.290 0.455 2.410 1.265 ;
        RECT  1.330 0.455 2.290 0.575 ;
        RECT  1.570 1.400 1.990 1.520 ;
        RECT  1.570 0.695 1.910 0.815 ;
        RECT  1.450 0.695 1.570 1.520 ;
        RECT  1.210 0.455 1.330 1.620 ;
        RECT  0.675 0.695 1.210 0.815 ;
        RECT  1.050 1.500 1.210 1.620 ;
    END
END AO2B2X1AD
MACRO AO2B2X2AD
    CLASS CORE ;
    FOREIGN AO2B2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.705 0.330 2.730 1.680 ;
        RECT  2.590 0.330 2.705 1.985 ;
        RECT  2.560 0.330 2.590 0.850 ;
        RECT  2.535 1.555 2.590 1.985 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 0.960 0.430 1.375 ;
        RECT  0.070 1.145 0.230 1.375 ;
        END
        AntennaGateArea 0.0834 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 0.960 0.770 1.375 ;
        END
        AntennaGateArea 0.0834 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.035 2.170 1.375 ;
        RECT  1.880 1.035 2.030 1.210 ;
        END
        AntennaGateArea 0.0603 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 0.960 1.090 1.375 ;
        END
        AntennaGateArea 0.0834 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.390 -0.210 2.800 0.210 ;
        RECT  2.130 -0.210 2.390 0.390 ;
        RECT  1.585 -0.210 2.130 0.210 ;
        RECT  1.325 -0.210 1.585 0.400 ;
        RECT  0.270 -0.210 1.325 0.210 ;
        RECT  0.100 -0.210 0.270 0.840 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.345 2.310 2.800 2.730 ;
        RECT  2.175 1.555 2.345 2.730 ;
        RECT  0.610 2.310 2.175 2.730 ;
        RECT  0.350 1.500 0.610 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.410 1.020 2.470 1.280 ;
        RECT  2.290 0.520 2.410 1.280 ;
        RECT  1.330 0.520 2.290 0.640 ;
        RECT  1.570 0.760 1.990 0.880 ;
        RECT  1.775 1.475 1.945 1.645 ;
        RECT  1.570 1.475 1.775 1.595 ;
        RECT  1.450 0.760 1.570 1.595 ;
        RECT  1.210 0.520 1.330 1.690 ;
        RECT  0.675 0.695 1.210 0.815 ;
        RECT  1.095 1.520 1.210 1.690 ;
    END
END AO2B2X2AD
MACRO AO2B2X4AD
    CLASS CORE ;
    FOREIGN AO2B2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.005 2.755 1.515 ;
        RECT  2.590 0.365 2.720 2.155 ;
        RECT  2.490 0.365 2.590 0.885 ;
        RECT  2.490 1.375 2.590 2.155 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.285 1.020 0.490 1.375 ;
        RECT  0.070 1.145 0.285 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.850 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.705 1.005 2.090 1.330 ;
        END
        AntennaGateArea 0.0674 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.980 0.865 1.330 1.275 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 -0.210 3.080 0.210 ;
        RECT  2.850 -0.210 2.970 0.865 ;
        RECT  2.320 -0.210 2.850 0.210 ;
        RECT  2.060 -0.210 2.320 0.390 ;
        RECT  1.620 -0.210 2.060 0.210 ;
        RECT  1.360 -0.210 1.620 0.390 ;
        RECT  0.325 -0.210 1.360 0.210 ;
        RECT  0.155 -0.210 0.325 0.785 ;
        RECT  0.000 -0.210 0.155 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 2.310 3.080 2.730 ;
        RECT  2.850 1.680 2.970 2.730 ;
        RECT  2.275 2.310 2.850 2.730 ;
        RECT  2.105 2.105 2.275 2.730 ;
        RECT  0.615 2.310 2.105 2.730 ;
        RECT  0.445 1.735 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  2.345 1.005 2.400 1.265 ;
        RECT  2.225 0.520 2.345 1.810 ;
        RECT  0.980 0.520 2.225 0.640 ;
        RECT  1.335 1.690 2.225 1.810 ;
        RECT  1.575 1.450 2.010 1.570 ;
        RECT  1.575 0.760 1.960 0.880 ;
        RECT  1.525 1.935 1.695 2.140 ;
        RECT  1.455 0.760 1.575 1.570 ;
        RECT  0.975 2.020 1.525 2.140 ;
        RECT  1.165 1.470 1.335 1.900 ;
        RECT  0.720 0.360 0.980 0.740 ;
        RECT  0.805 1.495 0.975 2.140 ;
        RECT  0.255 1.495 0.805 1.615 ;
        RECT  0.085 1.495 0.255 2.020 ;
    END
END AO2B2X4AD
MACRO AO2B2XLAD
    CLASS CORE ;
    FOREIGN AO2B2XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.670 2.730 1.650 ;
        RECT  2.535 0.670 2.590 0.840 ;
        RECT  2.535 1.480 2.590 1.650 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.395 1.280 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 0.865 0.770 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.865 2.170 1.245 ;
        RECT  1.915 0.975 2.030 1.245 ;
        END
        AntennaGateArea 0.0404 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 0.865 1.090 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.370 -0.210 2.800 0.210 ;
        RECT  2.110 -0.210 2.370 0.330 ;
        RECT  1.585 -0.210 2.110 0.210 ;
        RECT  1.325 -0.210 1.585 0.330 ;
        RECT  0.270 -0.210 1.325 0.210 ;
        RECT  0.100 -0.210 0.270 0.745 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.345 2.310 2.800 2.730 ;
        RECT  2.175 1.480 2.345 2.730 ;
        RECT  0.610 2.310 2.175 2.730 ;
        RECT  0.350 1.500 0.610 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.410 1.005 2.470 1.265 ;
        RECT  2.290 0.455 2.410 1.265 ;
        RECT  1.330 0.455 2.290 0.575 ;
        RECT  1.570 1.400 1.990 1.520 ;
        RECT  1.570 0.695 1.910 0.815 ;
        RECT  1.450 0.695 1.570 1.520 ;
        RECT  1.210 0.455 1.330 1.620 ;
        RECT  0.675 0.600 1.210 0.720 ;
        RECT  1.050 1.500 1.210 1.620 ;
    END
END AO2B2XLAD
MACRO AOI211X1AD
    CLASS CORE ;
    FOREIGN AOI211X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.535 1.585 0.870 ;
        RECT  1.415 1.495 1.585 1.925 ;
        RECT  1.290 0.750 1.415 0.870 ;
        RECT  1.330 1.495 1.415 1.655 ;
        RECT  1.290 1.425 1.330 1.655 ;
        RECT  1.170 0.750 1.290 1.655 ;
        RECT  0.865 0.750 1.170 0.870 ;
        RECT  0.695 0.535 0.865 0.870 ;
        END
        AntennaDiffArea 0.283 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 1.010 1.050 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 1.120 1.610 1.375 ;
        RECT  1.470 1.000 1.550 1.375 ;
        RECT  1.410 1.000 1.470 1.275 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.960 0.230 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.010 0.690 1.375 ;
        RECT  0.350 0.865 0.550 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.210 1.680 0.210 ;
        RECT  1.010 -0.210 1.270 0.630 ;
        RECT  0.255 -0.210 1.010 0.210 ;
        RECT  0.085 -0.210 0.255 0.710 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.660 2.310 1.680 2.730 ;
        RECT  0.400 1.760 0.660 2.730 ;
        RECT  0.000 2.310 0.400 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  0.805 1.495 0.975 1.955 ;
        RECT  0.255 1.495 0.805 1.615 ;
        RECT  0.085 1.495 0.255 1.925 ;
    END
END AOI211X1AD
MACRO AOI211X2AD
    CLASS CORE ;
    FOREIGN AOI211X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.460 1.585 0.745 ;
        RECT  1.350 1.520 1.560 2.040 ;
        RECT  1.290 0.625 1.415 0.745 ;
        RECT  1.290 1.425 1.350 2.040 ;
        RECT  1.170 0.625 1.290 2.040 ;
        RECT  0.910 0.625 1.170 0.745 ;
        RECT  0.650 0.365 0.910 0.745 ;
        END
        AntennaDiffArea 0.553 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.865 1.610 1.375 ;
        RECT  1.430 1.015 1.470 1.275 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.960 0.230 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.010 0.690 1.375 ;
        RECT  0.350 0.865 0.550 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 -0.210 1.680 0.210 ;
        RECT  1.055 -0.210 1.225 0.505 ;
        RECT  0.255 -0.210 1.055 0.210 ;
        RECT  0.085 -0.210 0.255 0.770 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.615 2.310 1.680 2.730 ;
        RECT  0.445 1.755 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  0.805 1.495 0.975 2.010 ;
        RECT  0.255 1.495 0.805 1.615 ;
        RECT  0.085 1.495 0.255 2.010 ;
    END
END AOI211X2AD
MACRO AOI211X4AD
    CLASS CORE ;
    FOREIGN AOI211X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.330 2.995 0.760 ;
        RECT  2.855 0.330 2.975 1.610 ;
        RECT  2.825 0.330 2.855 0.760 ;
        RECT  2.350 1.450 2.855 1.610 ;
        RECT  2.320 0.605 2.825 0.730 ;
        RECT  2.090 1.450 2.350 1.885 ;
        RECT  2.060 0.350 2.320 0.730 ;
        RECT  1.600 0.605 2.060 0.730 ;
        RECT  1.340 0.350 1.600 0.730 ;
        RECT  0.360 0.605 1.340 0.730 ;
        RECT  0.100 0.350 0.360 0.730 ;
        END
        AntennaDiffArea 0.92 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.615 0.850 2.735 1.280 ;
        RECT  1.890 0.850 2.615 0.970 ;
        RECT  1.640 0.850 1.890 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.140 1.110 2.495 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.090 1.130 1.355 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 0.850 1.440 1.280 ;
        RECT  0.490 0.850 1.320 0.970 ;
        RECT  0.210 0.850 0.490 1.275 ;
        RECT  0.070 0.850 0.210 1.095 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.635 -0.210 3.080 0.210 ;
        RECT  2.465 -0.210 2.635 0.465 ;
        RECT  1.915 -0.210 2.465 0.210 ;
        RECT  1.745 -0.210 1.915 0.460 ;
        RECT  0.970 -0.210 1.745 0.210 ;
        RECT  0.710 -0.210 0.970 0.485 ;
        RECT  0.000 -0.210 0.710 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.335 2.310 3.080 2.730 ;
        RECT  1.165 1.770 1.335 2.730 ;
        RECT  0.615 2.310 1.165 2.730 ;
        RECT  0.445 1.770 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  2.815 1.745 2.985 2.175 ;
        RECT  1.695 2.020 2.815 2.140 ;
        RECT  1.525 1.495 1.695 2.140 ;
        RECT  0.975 1.495 1.525 1.615 ;
        RECT  0.805 1.495 0.975 2.010 ;
        RECT  0.255 1.495 0.805 1.615 ;
        RECT  0.085 1.495 0.255 2.005 ;
    END
END AOI211X4AD
MACRO AOI211XLAD
    CLASS CORE ;
    FOREIGN AOI211XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.600 1.585 1.770 ;
        RECT  1.440 0.440 1.560 0.870 ;
        RECT  1.310 0.750 1.440 0.870 ;
        RECT  1.310 1.425 1.350 1.935 ;
        RECT  1.190 0.750 1.310 1.935 ;
        RECT  0.865 0.750 1.190 0.870 ;
        RECT  0.695 0.485 0.865 0.870 ;
        END
        AntennaDiffArea 0.193 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 1.010 1.050 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.570 1.130 1.610 1.475 ;
        RECT  1.470 0.995 1.570 1.475 ;
        RECT  1.430 0.995 1.470 1.275 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.830 0.230 1.375 ;
        END
        AntennaGateArea 0.062 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.010 0.690 1.375 ;
        RECT  0.350 0.865 0.550 1.375 ;
        END
        AntennaGateArea 0.062 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.210 1.680 0.210 ;
        RECT  1.010 -0.210 1.270 0.630 ;
        RECT  0.255 -0.210 1.010 0.210 ;
        RECT  0.085 -0.210 0.255 0.650 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.660 2.310 1.680 2.730 ;
        RECT  0.400 1.735 0.660 2.730 ;
        RECT  0.000 2.310 0.400 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  0.805 1.495 0.975 1.805 ;
        RECT  0.255 1.495 0.805 1.615 ;
        RECT  0.085 1.495 0.255 1.790 ;
    END
END AOI211XLAD
MACRO AOI21BX1AD
    CLASS CORE ;
    FOREIGN AOI21BX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.085 0.660 2.170 1.505 ;
        RECT  2.030 0.660 2.085 1.935 ;
        RECT  1.985 0.660 2.030 0.830 ;
        RECT  1.915 1.395 2.030 1.935 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.975 1.150 1.375 ;
        END
        AntennaGateArea 0.0414 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.055 0.225 1.655 ;
        END
        AntennaGateArea 0.0404 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.585 0.975 0.790 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.210 2.240 0.210 ;
        RECT  1.595 -0.210 1.765 0.505 ;
        RECT  0.905 -0.210 1.595 0.210 ;
        RECT  0.735 -0.210 0.905 0.420 ;
        RECT  0.000 -0.210 0.735 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 2.310 2.240 2.730 ;
        RECT  1.555 1.775 1.725 2.730 ;
        RECT  0.565 2.310 1.555 2.730 ;
        RECT  0.565 1.940 0.690 2.110 ;
        RECT  0.395 1.940 0.565 2.730 ;
        RECT  0.260 1.940 0.395 2.110 ;
        RECT  0.000 2.310 0.395 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.505 1.015 1.910 1.275 ;
        RECT  1.335 0.685 1.505 1.615 ;
        RECT  1.215 0.430 1.430 0.550 ;
        RECT  1.060 1.495 1.335 1.615 ;
        RECT  1.095 0.430 1.215 0.855 ;
        RECT  0.465 0.685 1.095 0.855 ;
        RECT  0.465 1.495 0.605 1.615 ;
        RECT  0.345 0.685 0.465 1.615 ;
        RECT  0.100 0.685 0.345 0.855 ;
    END
END AOI21BX1AD
MACRO AOI21BX2AD
    CLASS CORE ;
    FOREIGN AOI21BX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.345 2.170 2.140 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.015 1.160 1.375 ;
        END
        AntennaGateArea 0.0734 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.240 1.280 ;
        RECT  0.070 1.020 0.210 1.665 ;
        END
        AntennaGateArea 0.0604 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.015 0.790 1.380 ;
        END
        AntennaGateArea 0.0604 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.795 -0.210 2.240 0.210 ;
        RECT  1.625 -0.210 1.795 0.415 ;
        RECT  0.875 -0.210 1.625 0.210 ;
        RECT  0.705 -0.210 0.875 0.375 ;
        RECT  0.000 -0.210 0.705 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.705 2.310 2.240 2.730 ;
        RECT  1.535 1.755 1.705 2.730 ;
        RECT  0.895 2.310 1.535 2.730 ;
        RECT  0.725 1.925 0.895 2.730 ;
        RECT  0.255 2.310 0.725 2.730 ;
        RECT  0.085 1.925 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.515 1.015 1.870 1.275 ;
        RECT  1.345 0.655 1.515 1.620 ;
        RECT  1.215 0.330 1.440 0.450 ;
        RECT  1.060 1.500 1.345 1.620 ;
        RECT  1.095 0.330 1.215 0.880 ;
        RECT  0.480 0.760 1.095 0.880 ;
        RECT  0.480 1.500 0.620 1.620 ;
        RECT  0.360 0.760 0.480 1.620 ;
        RECT  0.270 0.760 0.360 0.880 ;
        RECT  0.100 0.710 0.270 0.880 ;
    END
END AOI21BX2AD
MACRO AOI21BX4AD
    CLASS CORE ;
    FOREIGN AOI21BX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.075 1.005 2.170 1.515 ;
        RECT  1.905 0.395 2.075 2.120 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 0.585 1.050 1.240 ;
        END
        AntennaGateArea 0.1444 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.235 1.015 0.380 1.275 ;
        RECT  0.210 1.145 0.235 1.275 ;
        RECT  0.070 1.145 0.210 1.375 ;
        END
        AntennaGateArea 0.0684 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.495 1.705 0.770 2.050 ;
        END
        AntennaGateArea 0.0684 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 -0.210 2.520 0.210 ;
        RECT  2.265 -0.210 2.435 0.830 ;
        RECT  1.715 -0.210 2.265 0.210 ;
        RECT  1.545 -0.210 1.715 0.480 ;
        RECT  0.765 -0.210 1.545 0.210 ;
        RECT  0.595 -0.210 0.765 0.345 ;
        RECT  0.000 -0.210 0.595 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 2.310 2.520 2.730 ;
        RECT  2.265 1.625 2.435 2.730 ;
        RECT  1.635 2.310 2.265 2.730 ;
        RECT  1.465 1.865 1.635 2.730 ;
        RECT  0.870 2.310 1.465 2.730 ;
        RECT  0.610 2.175 0.870 2.730 ;
        RECT  0.255 2.310 0.610 2.730 ;
        RECT  0.085 1.955 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.640 0.695 1.760 1.730 ;
        RECT  1.275 0.695 1.640 0.865 ;
        RECT  1.215 1.610 1.640 1.730 ;
        RECT  1.220 1.000 1.340 1.490 ;
        RECT  0.620 1.370 1.220 1.490 ;
        RECT  1.045 1.610 1.215 2.040 ;
        RECT  0.500 0.765 0.620 1.585 ;
        RECT  0.255 0.765 0.500 0.885 ;
        RECT  0.375 1.415 0.500 1.585 ;
        RECT  0.085 0.685 0.255 0.885 ;
    END
END AOI21BX4AD
MACRO AOI21BXLAD
    CLASS CORE ;
    FOREIGN AOI21BXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.610 2.170 1.785 ;
        RECT  1.975 0.610 2.030 0.780 ;
        RECT  1.915 1.615 2.030 1.785 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.900 0.975 1.150 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.055 0.225 1.655 ;
        END
        AntennaGateArea 0.0404 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.585 0.975 0.775 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.755 -0.210 2.240 0.210 ;
        RECT  1.585 -0.210 1.755 0.505 ;
        RECT  0.905 -0.210 1.585 0.210 ;
        RECT  0.735 -0.210 0.905 0.420 ;
        RECT  0.000 -0.210 0.735 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.675 2.310 2.240 2.730 ;
        RECT  1.675 1.735 1.740 1.855 ;
        RECT  1.535 1.735 1.675 2.730 ;
        RECT  1.480 1.735 1.535 1.855 ;
        RECT  0.565 2.310 1.535 2.730 ;
        RECT  0.565 1.940 0.690 2.110 ;
        RECT  0.395 1.940 0.565 2.730 ;
        RECT  0.260 1.940 0.395 2.110 ;
        RECT  0.000 2.310 0.395 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.790 0.895 1.910 1.415 ;
        RECT  1.505 1.095 1.790 1.255 ;
        RECT  1.335 0.685 1.505 1.615 ;
        RECT  1.215 0.430 1.430 0.550 ;
        RECT  1.320 1.495 1.335 1.615 ;
        RECT  1.060 1.495 1.320 1.655 ;
        RECT  1.095 0.430 1.215 0.855 ;
        RECT  0.465 0.685 1.095 0.855 ;
        RECT  0.465 1.535 0.605 1.655 ;
        RECT  0.345 0.685 0.465 1.655 ;
        RECT  0.100 0.685 0.345 0.855 ;
    END
END AOI21BXLAD
MACRO AOI21X1AD
    CLASS CORE ;
    FOREIGN AOI21X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.625 1.330 1.925 ;
        RECT  0.670 0.625 1.170 0.745 ;
        END
        AntennaDiffArea 0.222 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 1.020 1.050 1.655 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.405 1.230 ;
        RECT  0.070 1.020 0.210 1.655 ;
        END
        AntennaGateArea 0.0884 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 0.865 0.770 1.375 ;
        END
        AntennaGateArea 0.0904 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.295 -0.210 1.400 0.210 ;
        RECT  1.125 -0.210 1.295 0.505 ;
        RECT  0.275 -0.210 1.125 0.210 ;
        RECT  0.105 -0.210 0.275 0.820 ;
        RECT  0.000 -0.210 0.105 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.310 1.400 2.730 ;
        RECT  0.360 2.230 0.620 2.730 ;
        RECT  0.000 2.310 0.360 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.105 1.775 1.000 1.945 ;
    END
END AOI21X1AD
MACRO AOI21X2AD
    CLASS CORE ;
    FOREIGN AOI21X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.785 1.610 1.655 ;
        RECT  0.915 0.785 1.470 0.905 ;
        RECT  1.375 1.535 1.470 1.655 ;
        RECT  1.205 1.535 1.375 1.990 ;
        RECT  0.745 0.400 0.915 0.905 ;
        END
        AntennaDiffArea 0.408 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.040 1.330 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.270 1.020 0.440 1.375 ;
        RECT  0.070 1.145 0.270 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 1.025 0.780 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.395 -0.210 1.680 0.210 ;
        RECT  1.395 0.475 1.545 0.645 ;
        RECT  1.240 -0.210 1.395 0.645 ;
        RECT  0.295 -0.210 1.240 0.210 ;
        RECT  1.115 0.475 1.240 0.645 ;
        RECT  0.125 -0.210 0.295 0.815 ;
        RECT  0.000 -0.210 0.125 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.655 2.310 1.680 2.730 ;
        RECT  0.485 1.735 0.655 2.730 ;
        RECT  0.000 2.310 0.485 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  0.845 1.495 1.015 2.005 ;
        RECT  0.305 1.495 0.845 1.615 ;
        RECT  0.125 1.495 0.305 2.035 ;
    END
END AOI21X2AD
MACRO AOI21X3AD
    CLASS CORE ;
    FOREIGN AOI21X3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.410 0.770 2.450 1.615 ;
        RECT  2.310 0.565 2.410 1.615 ;
        RECT  2.230 0.565 2.310 0.890 ;
        RECT  2.120 1.495 2.310 1.615 ;
        RECT  1.640 0.770 2.230 0.890 ;
        RECT  1.860 1.495 2.120 1.875 ;
        RECT  1.470 0.600 1.640 0.890 ;
        RECT  0.315 0.770 1.470 0.890 ;
        RECT  0.145 0.610 0.315 0.890 ;
        END
        AntennaDiffArea 0.62 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.045 2.190 1.375 ;
        END
        AntennaGateArea 0.244 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.065 1.105 1.330 ;
        END
        AntennaGateArea 0.244 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.305 1.045 1.475 1.570 ;
        RECT  0.530 1.450 1.305 1.570 ;
        RECT  0.390 1.035 0.530 1.570 ;
        RECT  0.320 1.035 0.390 1.375 ;
        RECT  0.070 1.145 0.320 1.375 ;
        END
        AntennaGateArea 0.244 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.075 -0.210 2.520 0.210 ;
        RECT  1.905 -0.210 2.075 0.650 ;
        RECT  0.955 -0.210 1.905 0.210 ;
        RECT  0.785 -0.210 0.955 0.650 ;
        RECT  0.000 -0.210 0.785 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 2.310 2.520 2.730 ;
        RECT  1.330 1.930 1.400 2.050 ;
        RECT  1.210 1.930 1.330 2.730 ;
        RECT  1.140 1.930 1.210 2.050 ;
        RECT  0.600 2.310 1.210 2.730 ;
        RECT  0.600 1.930 0.670 2.050 ;
        RECT  0.480 1.930 0.600 2.730 ;
        RECT  0.410 1.930 0.480 2.050 ;
        RECT  0.000 2.310 0.480 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.265 1.735 2.435 2.115 ;
        RECT  1.715 1.995 2.265 2.115 ;
        RECT  1.545 1.690 1.715 2.115 ;
        RECT  0.230 1.690 1.545 1.810 ;
        RECT  0.110 1.500 0.230 2.020 ;
    END
END AOI21X3AD
MACRO AOI21X4AD
    CLASS CORE ;
    FOREIGN AOI21X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.410 0.630 2.450 1.545 ;
        RECT  2.290 0.330 2.410 1.545 ;
        RECT  1.610 0.630 2.290 0.760 ;
        RECT  2.055 1.405 2.290 1.545 ;
        RECT  1.885 1.405 2.055 1.880 ;
        RECT  1.440 0.330 1.610 0.760 ;
        RECT  0.365 0.630 1.440 0.760 ;
        RECT  0.195 0.330 0.365 0.760 ;
        END
        AntennaDiffArea 0.802 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.705 0.910 2.170 1.230 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.120 1.160 1.240 ;
        RECT  0.630 1.120 1.050 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.335 0.880 1.455 1.260 ;
        RECT  0.490 0.880 1.335 1.000 ;
        RECT  0.295 0.880 0.490 1.375 ;
        RECT  0.070 1.145 0.295 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.055 -0.210 2.520 0.210 ;
        RECT  1.885 -0.210 2.055 0.505 ;
        RECT  0.985 -0.210 1.885 0.210 ;
        RECT  0.815 -0.210 0.985 0.510 ;
        RECT  0.000 -0.210 0.815 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.335 2.310 2.520 2.730 ;
        RECT  1.165 1.845 1.335 2.730 ;
        RECT  0.615 2.310 1.165 2.730 ;
        RECT  0.445 1.795 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.265 1.710 2.435 2.140 ;
        RECT  1.695 2.020 2.265 2.140 ;
        RECT  1.525 1.520 1.695 2.140 ;
        RECT  0.975 1.520 1.525 1.640 ;
        RECT  0.805 1.520 0.975 1.980 ;
        RECT  0.255 1.520 0.805 1.640 ;
        RECT  0.085 1.520 0.255 1.980 ;
    END
END AOI21X4AD
MACRO AOI21X6AD
    CLASS CORE ;
    FOREIGN AOI21X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.495 0.805 3.570 1.655 ;
        RECT  3.400 0.805 3.495 2.140 ;
        RECT  3.385 0.805 3.400 0.985 ;
        RECT  3.295 1.515 3.400 2.140 ;
        RECT  3.215 0.410 3.385 0.985 ;
        RECT  2.820 1.960 3.295 2.140 ;
        RECT  2.665 0.805 3.215 0.985 ;
        RECT  2.560 1.760 2.820 2.140 ;
        RECT  2.495 0.425 2.665 0.985 ;
        RECT  1.670 0.620 2.495 0.780 ;
        RECT  1.410 0.400 1.670 0.780 ;
        RECT  0.365 0.620 1.410 0.780 ;
        RECT  0.195 0.420 0.365 0.850 ;
        END
        AntennaDiffArea 1.21 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 1.120 3.150 1.240 ;
        RECT  2.590 1.120 3.010 1.375 ;
        RECT  2.370 1.120 2.590 1.240 ;
        END
        AntennaGateArea 0.486 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.985 0.900 2.155 1.250 ;
        RECT  1.120 0.900 1.985 1.020 ;
        RECT  0.715 0.900 1.120 1.330 ;
        END
        AntennaGateArea 0.486 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.410 1.140 1.825 1.260 ;
        RECT  1.285 1.140 1.410 1.570 ;
        RECT  0.490 1.450 1.285 1.570 ;
        RECT  0.325 1.015 0.490 1.570 ;
        RECT  0.260 1.145 0.325 1.570 ;
        RECT  0.070 1.145 0.260 1.375 ;
        END
        AntennaGateArea 0.4869 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.025 -0.210 3.640 0.210 ;
        RECT  2.855 -0.210 3.025 0.675 ;
        RECT  2.350 -0.210 2.855 0.210 ;
        RECT  2.090 -0.210 2.350 0.500 ;
        RECT  1.020 -0.210 2.090 0.210 ;
        RECT  0.760 -0.210 1.020 0.500 ;
        RECT  0.000 -0.210 0.760 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.055 2.310 3.640 2.730 ;
        RECT  1.885 1.735 2.055 2.730 ;
        RECT  1.335 2.310 1.885 2.730 ;
        RECT  1.165 1.930 1.335 2.730 ;
        RECT  0.615 2.310 1.165 2.730 ;
        RECT  0.445 1.930 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  2.965 1.495 3.135 1.835 ;
        RECT  2.415 1.495 2.965 1.615 ;
        RECT  2.245 1.495 2.415 2.010 ;
        RECT  1.695 1.495 2.245 1.615 ;
        RECT  1.565 1.495 1.695 2.120 ;
        RECT  1.525 1.690 1.565 2.120 ;
        RECT  0.975 1.690 1.525 1.810 ;
        RECT  0.805 1.690 0.975 2.120 ;
        RECT  0.255 1.690 0.805 1.810 ;
        RECT  0.085 1.690 0.255 2.120 ;
    END
END AOI21X6AD
MACRO AOI21X8AD
    CLASS CORE ;
    FOREIGN AOI21X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.280 0.800 4.550 1.760 ;
        RECT  4.260 0.370 4.280 1.760 ;
        RECT  4.130 0.370 4.260 1.875 ;
        RECT  4.050 0.370 4.130 0.960 ;
        RECT  4.000 1.495 4.130 1.875 ;
        RECT  3.505 0.620 4.050 0.960 ;
        RECT  3.540 1.495 4.000 1.760 ;
        RECT  3.280 1.495 3.540 1.875 ;
        RECT  3.280 0.380 3.505 0.960 ;
        RECT  2.470 0.620 3.280 0.780 ;
        RECT  2.210 0.400 2.470 0.780 ;
        RECT  1.030 0.620 2.210 0.780 ;
        RECT  0.770 0.400 1.030 0.780 ;
        END
        AntennaDiffArea 1.236 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.595 1.135 3.940 1.255 ;
        RECT  3.150 1.135 3.595 1.375 ;
        END
        AntennaGateArea 0.6499 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.755 0.900 2.925 1.255 ;
        RECT  1.810 0.900 2.755 1.020 ;
        RECT  1.425 0.900 1.810 1.330 ;
        RECT  0.465 0.900 1.425 1.020 ;
        RECT  0.295 0.900 0.465 1.275 ;
        END
        AntennaGateArea 0.648 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.125 1.140 2.600 1.260 ;
        RECT  2.000 1.140 2.125 1.570 ;
        RECT  1.050 1.450 2.000 1.570 ;
        RECT  0.930 1.140 1.050 1.570 ;
        RECT  0.630 1.140 0.930 1.375 ;
        END
        AntennaGateArea 0.6499 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.580 -0.210 4.760 0.210 ;
        RECT  4.410 -0.210 4.580 0.675 ;
        RECT  3.860 -0.210 4.410 0.210 ;
        RECT  3.690 -0.210 3.860 0.490 ;
        RECT  3.125 -0.210 3.690 0.210 ;
        RECT  2.865 -0.210 3.125 0.500 ;
        RECT  1.775 -0.210 2.865 0.210 ;
        RECT  1.465 -0.210 1.775 0.500 ;
        RECT  0.365 -0.210 1.465 0.210 ;
        RECT  0.195 -0.210 0.365 0.775 ;
        RECT  0.000 -0.210 0.195 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.775 2.310 4.760 2.730 ;
        RECT  2.605 1.735 2.775 2.730 ;
        RECT  2.055 2.310 2.605 2.730 ;
        RECT  1.885 1.930 2.055 2.730 ;
        RECT  1.335 2.310 1.885 2.730 ;
        RECT  1.165 1.930 1.335 2.730 ;
        RECT  0.615 2.310 1.165 2.730 ;
        RECT  0.445 1.950 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.760 2.520 ;
        LAYER M1 ;
        RECT  4.410 1.885 4.580 2.140 ;
        RECT  3.135 2.020 4.410 2.140 ;
        RECT  2.965 1.495 3.135 2.185 ;
        RECT  2.415 1.495 2.965 1.615 ;
        RECT  2.245 1.495 2.415 2.045 ;
        RECT  1.695 1.690 2.245 1.810 ;
        RECT  1.525 1.690 1.695 2.120 ;
        RECT  1.020 1.690 1.525 1.810 ;
        RECT  0.760 1.690 1.020 2.070 ;
        RECT  0.255 1.690 0.760 1.810 ;
        RECT  0.085 1.415 0.255 2.105 ;
    END
END AOI21X8AD
MACRO AOI21XLAD
    CLASS CORE ;
    FOREIGN AOI21XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.780 1.330 1.715 ;
        RECT  0.885 0.780 1.170 0.900 ;
        RECT  0.715 0.730 0.885 0.900 ;
        END
        AntennaDiffArea 0.156 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.020 1.050 1.655 ;
        END
        AntennaGateArea 0.0604 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.400 1.280 ;
        RECT  0.130 1.020 0.210 1.655 ;
        RECT  0.070 1.145 0.130 1.655 ;
        END
        AntennaGateArea 0.0604 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 1.020 0.770 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.270 -0.210 1.400 0.210 ;
        RECT  1.100 -0.210 1.270 0.660 ;
        RECT  0.270 -0.210 1.100 0.210 ;
        RECT  0.100 -0.210 0.270 0.900 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.575 2.310 1.400 2.730 ;
        RECT  0.405 1.515 0.575 2.730 ;
        RECT  0.000 2.310 0.405 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
	 END
END AOI21XLAD
MACRO AOI221X1AD
    CLASS CORE ;
    FOREIGN AOI221X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.435 0.780 2.450 1.605 ;
        RECT  2.365 0.780 2.435 1.925 ;
        RECT  2.310 0.560 2.365 1.925 ;
        RECT  2.195 0.560 2.310 0.900 ;
        RECT  2.265 1.495 2.310 1.925 ;
        RECT  1.635 0.780 2.195 0.900 ;
        RECT  1.515 0.585 1.635 0.900 ;
        RECT  0.825 0.585 1.515 0.705 ;
        END
        AntennaDiffArea 0.387 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.020 2.190 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.965 0.465 1.225 ;
        RECT  0.240 0.965 0.350 1.375 ;
        RECT  0.070 1.145 0.240 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.585 0.910 0.885 1.240 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.020 1.890 1.395 ;
        RECT  1.645 1.020 1.750 1.240 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.145 0.910 1.395 1.240 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.020 -0.210 2.520 0.210 ;
        RECT  1.760 -0.210 2.020 0.660 ;
        RECT  0.395 -0.210 1.760 0.210 ;
        RECT  0.225 -0.210 0.395 0.730 ;
        RECT  0.000 -0.210 0.225 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.005 2.310 2.520 2.730 ;
        RECT  0.835 1.600 1.005 2.730 ;
        RECT  0.280 2.310 0.835 2.730 ;
        RECT  0.110 1.525 0.280 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.905 1.525 2.075 1.955 ;
        RECT  1.345 1.835 1.905 1.955 ;
        RECT  1.630 1.535 1.715 1.705 ;
        RECT  1.510 1.360 1.630 1.705 ;
        RECT  0.645 1.360 1.510 1.480 ;
        RECT  1.175 1.615 1.345 1.955 ;
        RECT  0.475 1.360 0.645 1.850 ;
    END
END AOI221X1AD
MACRO AOI221X2AD
    CLASS CORE ;
    FOREIGN AOI221X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.435 0.625 2.450 1.570 ;
        RECT  2.310 0.340 2.435 2.160 ;
        RECT  2.265 0.340 2.310 0.770 ;
        RECT  2.265 1.470 2.310 2.160 ;
        RECT  1.390 0.625 2.265 0.745 ;
        RECT  0.960 0.480 1.390 0.745 ;
        END
        AntennaDiffArea 0.869 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.865 2.190 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 1.010 0.440 1.375 ;
        RECT  0.070 1.120 0.295 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.585 0.910 0.900 1.330 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.865 1.910 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.145 0.910 1.585 1.330 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.075 -0.210 2.520 0.210 ;
        RECT  1.905 -0.210 2.075 0.505 ;
        RECT  0.395 -0.210 1.905 0.210 ;
        RECT  0.225 -0.210 0.395 0.815 ;
        RECT  0.000 -0.210 0.225 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.005 2.310 2.520 2.730 ;
        RECT  0.835 1.760 1.005 2.730 ;
        RECT  0.285 2.310 0.835 2.730 ;
        RECT  0.115 1.525 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.905 1.595 2.075 2.140 ;
        RECT  1.345 2.020 1.905 2.140 ;
        RECT  1.500 1.510 1.760 1.890 ;
        RECT  0.645 1.510 1.500 1.630 ;
        RECT  1.175 1.750 1.345 2.180 ;
        RECT  0.475 1.510 0.645 2.015 ;
    END
END AOI221X2AD
MACRO AOI221X4AD
    CLASS CORE ;
    FOREIGN AOI221X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.035 0.660 4.130 1.900 ;
        RECT  3.990 0.360 4.035 1.900 ;
        RECT  3.865 0.360 3.990 0.790 ;
        RECT  3.820 1.520 3.990 1.900 ;
        RECT  2.955 0.660 3.865 0.790 ;
        RECT  2.785 0.360 2.955 0.790 ;
        RECT  1.640 0.660 2.785 0.790 ;
        RECT  1.520 0.385 1.640 0.790 ;
        RECT  0.770 0.385 1.520 0.505 ;
        END
        AntennaDiffArea 0.81 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.595 1.030 3.860 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.400 0.980 1.460 1.240 ;
        RECT  1.280 0.625 1.400 1.240 ;
        RECT  0.490 0.625 1.280 0.745 ;
        RECT  0.350 0.625 0.490 1.250 ;
        RECT  0.070 0.865 0.350 1.095 ;
        END
        AntennaGateArea 0.324 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.050 1.160 1.170 ;
        RECT  0.630 0.865 1.050 1.170 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.315 1.040 3.435 1.425 ;
        RECT  3.105 1.190 3.315 1.425 ;
        RECT  2.455 1.305 3.105 1.425 ;
        RECT  2.335 1.040 2.455 1.425 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.925 0.910 3.055 1.050 ;
        RECT  2.665 0.910 2.925 1.170 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.370 -0.210 4.480 0.210 ;
        RECT  4.250 -0.210 4.370 0.830 ;
        RECT  3.630 -0.210 4.250 0.210 ;
        RECT  3.460 -0.210 3.630 0.535 ;
        RECT  2.085 -0.210 3.460 0.210 ;
        RECT  2.085 0.370 2.190 0.540 ;
        RECT  1.895 -0.210 2.085 0.540 ;
        RECT  0.410 -0.210 1.895 0.210 ;
        RECT  1.760 0.370 1.895 0.540 ;
        RECT  0.150 -0.210 0.410 0.505 ;
        RECT  0.000 -0.210 0.150 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.695 2.310 4.480 2.730 ;
        RECT  1.525 1.660 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.725 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.465 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
        LAYER M1 ;
        RECT  4.250 1.555 4.370 2.140 ;
        RECT  3.675 2.020 4.250 2.140 ;
        RECT  3.505 1.615 3.675 2.140 ;
        RECT  2.065 1.970 3.505 2.140 ;
        RECT  2.215 1.610 3.315 1.780 ;
        RECT  2.095 1.415 2.215 1.780 ;
        RECT  1.335 1.415 2.095 1.535 ;
        RECT  1.165 1.415 1.335 1.975 ;
        RECT  0.615 1.415 1.165 1.535 ;
        RECT  0.445 1.415 0.615 1.990 ;
    END
END AOI221X4AD
MACRO AOI221XLAD
    CLASS CORE ;
    FOREIGN AOI221XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.155 0.555 2.170 1.935 ;
        RECT  2.050 0.505 2.155 1.935 ;
        RECT  1.985 0.505 2.050 0.675 ;
        RECT  2.030 1.425 2.050 1.935 ;
        RECT  1.985 1.535 2.030 1.705 ;
        RECT  0.975 0.555 1.985 0.675 ;
        RECT  0.805 0.505 0.975 0.675 ;
        END
        AntennaDiffArea 0.236 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 0.795 1.920 1.315 ;
        RECT  1.750 0.795 1.890 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.795 0.370 1.330 ;
        RECT  0.210 1.140 0.250 1.330 ;
        RECT  0.070 1.140 0.210 1.655 ;
        END
        AntennaGateArea 0.0604 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.795 0.770 1.375 ;
        RECT  0.580 0.795 0.630 1.315 ;
        END
        AntennaGateArea 0.0604 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.795 1.610 1.375 ;
        RECT  1.420 0.795 1.470 1.315 ;
        END
        AntennaGateArea 0.0604 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.795 1.230 1.315 ;
        RECT  0.910 0.795 1.050 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.800 -0.210 2.240 0.210 ;
        RECT  1.540 -0.210 1.800 0.435 ;
        RECT  0.265 -0.210 1.540 0.210 ;
        RECT  0.095 -0.210 0.265 0.675 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.570 2.310 2.240 2.730 ;
        RECT  0.570 2.065 0.870 2.185 ;
        RECT  0.350 2.065 0.570 2.730 ;
        RECT  0.090 2.065 0.350 2.185 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  0.375 1.535 1.475 1.705 ;
    END
END AOI221XLAD
MACRO AOI222X1AD
    CLASS CORE ;
    FOREIGN AOI222X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.700 2.730 1.635 ;
        RECT  1.985 0.700 2.590 0.820 ;
        RECT  2.400 1.495 2.590 1.635 ;
        RECT  2.140 1.495 2.400 1.875 ;
        RECT  1.765 0.625 1.985 0.820 ;
        RECT  0.255 0.625 1.765 0.745 ;
        RECT  0.085 0.625 0.255 0.840 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.545 0.865 0.770 1.250 ;
        END
        AntennaGateArea 0.09 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.970 0.380 1.250 ;
        RECT  0.115 0.970 0.210 1.375 ;
        RECT  0.070 1.130 0.115 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.865 1.350 1.250 ;
        END
        AntennaGateArea 0.09 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.645 0.990 1.760 1.250 ;
        RECT  1.470 0.865 1.645 1.250 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.940 2.470 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.915 0.940 2.170 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.670 -0.210 2.800 0.210 ;
        RECT  2.410 -0.210 2.670 0.580 ;
        RECT  1.070 -0.210 2.410 0.210 ;
        RECT  1.070 0.360 1.245 0.480 ;
        RECT  0.905 -0.210 1.070 0.480 ;
        RECT  0.000 -0.210 0.905 0.210 ;
        RECT  0.725 0.360 0.905 0.480 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.975 2.310 2.800 2.730 ;
        RECT  0.805 1.885 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.600 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.545 1.785 2.715 2.115 ;
        RECT  1.995 1.995 2.545 2.115 ;
        RECT  1.825 1.500 1.995 2.115 ;
        RECT  1.320 1.995 1.825 2.115 ;
        RECT  1.465 1.370 1.635 1.855 ;
        RECT  0.615 1.370 1.465 1.490 ;
        RECT  1.200 1.610 1.320 2.115 ;
        RECT  1.060 1.610 1.200 1.730 ;
        RECT  0.445 1.370 0.615 1.950 ;
    END
END AOI222X1AD
MACRO AOI222X2AD
    CLASS CORE ;
    FOREIGN AOI222X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.770 2.730 1.665 ;
        RECT  1.945 0.770 2.590 0.890 ;
        RECT  2.400 1.495 2.590 1.665 ;
        RECT  2.380 1.495 2.400 1.900 ;
        RECT  2.140 1.520 2.380 1.900 ;
        RECT  1.775 0.340 1.945 0.890 ;
        RECT  0.365 0.625 1.775 0.745 ;
        RECT  0.195 0.405 0.365 0.835 ;
        END
        AntennaDiffArea 0.649 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.960 1.260 ;
        END
        AntennaGateArea 0.162 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.000 0.470 1.260 ;
        RECT  0.070 1.000 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 0.865 1.350 1.250 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.070 1.800 1.190 ;
        RECT  1.470 0.865 1.610 1.190 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 1.020 2.470 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 1.065 2.170 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.640 -0.210 2.800 0.210 ;
        RECT  2.380 -0.210 2.640 0.650 ;
        RECT  1.110 -0.210 2.380 0.210 ;
        RECT  1.110 0.380 1.290 0.500 ;
        RECT  0.915 -0.210 1.110 0.500 ;
        RECT  0.000 -0.210 0.915 0.210 ;
        RECT  0.770 0.380 0.915 0.500 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.975 2.310 2.800 2.730 ;
        RECT  0.805 1.985 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.610 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.545 1.810 2.715 2.140 ;
        RECT  1.995 2.020 2.545 2.140 ;
        RECT  1.825 1.615 1.995 2.140 ;
        RECT  1.275 2.020 1.825 2.140 ;
        RECT  1.465 1.380 1.635 1.835 ;
        RECT  0.615 1.380 1.465 1.500 ;
        RECT  1.105 1.620 1.275 2.140 ;
        RECT  0.445 1.380 0.615 1.935 ;
    END
END AOI222X2AD
MACRO AOI222X4AD
    CLASS CORE ;
    FOREIGN AOI222X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.830 0.660 4.970 1.685 ;
        RECT  4.235 0.660 4.830 0.790 ;
        RECT  4.640 1.505 4.830 1.685 ;
        RECT  4.380 1.505 4.640 1.885 ;
        RECT  3.920 1.505 4.380 1.685 ;
        RECT  4.065 0.360 4.235 0.790 ;
        RECT  2.810 0.660 4.065 0.790 ;
        RECT  3.660 1.505 3.920 1.885 ;
        RECT  2.640 0.360 2.810 0.790 ;
        RECT  1.625 0.660 2.640 0.790 ;
        RECT  1.495 0.380 1.625 0.790 ;
        RECT  0.760 0.380 1.495 0.500 ;
        END
        AntennaDiffArea 1.038 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.070 1.510 1.190 ;
        RECT  1.250 0.620 1.370 1.190 ;
        RECT  0.490 0.620 1.250 0.740 ;
        RECT  0.350 0.620 0.490 1.240 ;
        RECT  0.295 0.865 0.350 1.240 ;
        RECT  0.070 0.865 0.295 1.095 ;
        END
        AntennaGateArea 0.324 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.050 1.130 1.170 ;
        RECT  0.610 0.865 1.050 1.170 ;
        END
        AntennaGateArea 0.324 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.130 1.035 3.275 1.400 ;
        RECT  2.285 1.280 3.130 1.400 ;
        RECT  2.035 0.910 2.285 1.400 ;
        RECT  1.705 0.910 2.035 1.050 ;
        END
        AntennaGateArea 0.324 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.855 1.040 2.980 1.160 ;
        RECT  2.525 0.910 2.855 1.160 ;
        RECT  2.460 1.040 2.525 1.160 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.435 1.040 4.670 1.380 ;
        RECT  3.730 1.260 4.435 1.380 ;
        RECT  3.430 1.040 3.730 1.380 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.945 0.910 4.290 1.140 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.845 -0.210 5.040 0.210 ;
        RECT  4.675 -0.210 4.845 0.540 ;
        RECT  3.605 -0.210 4.675 0.210 ;
        RECT  3.340 -0.210 3.605 0.510 ;
        RECT  2.065 -0.210 3.340 0.210 ;
        RECT  1.800 -0.210 2.065 0.540 ;
        RECT  0.410 -0.210 1.800 0.210 ;
        RECT  0.150 -0.210 0.410 0.500 ;
        RECT  0.000 -0.210 0.150 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.695 2.310 5.040 2.730 ;
        RECT  1.525 1.735 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.610 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.560 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.040 2.520 ;
        LAYER M1 ;
        RECT  4.785 1.835 4.955 2.140 ;
        RECT  4.235 2.005 4.785 2.140 ;
        RECT  4.065 1.845 4.235 2.140 ;
        RECT  3.515 2.005 4.065 2.140 ;
        RECT  3.345 1.595 3.515 2.140 ;
        RECT  2.795 2.020 3.345 2.140 ;
        RECT  2.940 1.520 3.200 1.900 ;
        RECT  2.480 1.520 2.940 1.640 ;
        RECT  2.625 1.760 2.795 2.190 ;
        RECT  2.075 2.020 2.625 2.140 ;
        RECT  2.220 1.520 2.480 1.900 ;
        RECT  1.910 1.520 2.220 1.640 ;
        RECT  1.905 1.760 2.075 2.190 ;
        RECT  1.790 1.360 1.910 1.640 ;
        RECT  1.335 1.360 1.790 1.480 ;
        RECT  1.165 1.360 1.335 2.015 ;
        RECT  0.615 1.360 1.165 1.480 ;
        RECT  0.445 1.360 0.615 2.015 ;
    END
END AOI222X4AD
MACRO AOI222XLAD
    CLASS CORE ;
    FOREIGN AOI222XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 0.625 2.450 1.935 ;
        RECT  0.270 0.625 2.330 0.745 ;
        RECT  2.310 1.425 2.330 1.935 ;
        RECT  1.965 1.510 2.310 1.680 ;
        RECT  0.100 0.600 0.270 0.770 ;
        END
        AntennaDiffArea 0.214 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.565 0.865 0.770 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.975 0.370 1.265 ;
        RECT  0.205 0.975 0.210 1.655 ;
        RECT  0.070 1.115 0.205 1.655 ;
        END
        AntennaGateArea 0.0604 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.865 1.070 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.050 1.610 1.170 ;
        RECT  1.190 0.865 1.330 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.200 0.925 2.210 1.185 ;
        RECT  2.175 0.865 2.200 1.185 ;
        RECT  2.030 0.865 2.175 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 0.865 1.900 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.405 -0.210 2.520 0.210 ;
        RECT  2.235 -0.210 2.405 0.505 ;
        RECT  1.035 -0.210 2.235 0.210 ;
        RECT  0.775 -0.210 1.035 0.505 ;
        RECT  0.000 -0.210 0.775 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.575 2.310 2.520 2.730 ;
        RECT  0.575 2.040 0.870 2.160 ;
        RECT  0.365 2.040 0.575 2.730 ;
        RECT  0.090 2.040 0.365 2.160 ;
        RECT  0.000 2.310 0.365 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  0.375 1.495 1.465 1.665 ;
    END
END AOI222XLAD
MACRO AOI22X1AD
    CLASS CORE ;
    FOREIGN AOI22X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.625 1.890 1.615 ;
        RECT  1.010 0.625 1.750 0.745 ;
        RECT  1.490 1.495 1.750 1.615 ;
        RECT  1.230 1.495 1.490 1.875 ;
        RECT  0.840 0.575 1.010 0.745 ;
        END
        AntennaDiffArea 0.266 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.000 0.485 1.260 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.605 0.865 0.790 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.385 0.865 1.610 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.865 1.210 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.715 -0.210 1.960 0.210 ;
        RECT  1.545 -0.210 1.715 0.500 ;
        RECT  0.360 -0.210 1.545 0.210 ;
        RECT  0.190 -0.210 0.360 0.740 ;
        RECT  0.000 -0.210 0.190 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.725 2.310 1.960 2.730 ;
        RECT  0.555 1.745 0.725 2.730 ;
        RECT  0.000 2.310 0.555 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.635 1.735 1.805 2.115 ;
        RECT  1.085 1.995 1.635 2.115 ;
        RECT  0.915 1.495 1.085 2.115 ;
        RECT  0.360 1.495 0.915 1.615 ;
        RECT  0.190 1.495 0.360 1.925 ;
    END
END AOI22X1AD
MACRO AOI22X2AD
    CLASS CORE ;
    FOREIGN AOI22X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.625 1.890 1.615 ;
        RECT  1.055 0.625 1.750 0.745 ;
        RECT  1.490 1.495 1.750 1.615 ;
        RECT  1.230 1.495 1.490 1.875 ;
        RECT  0.795 0.365 1.055 0.745 ;
        END
        AntennaDiffArea 0.5 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.045 0.465 1.215 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.865 0.790 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 0.865 1.610 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.865 1.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.695 -0.210 1.960 0.210 ;
        RECT  1.525 -0.210 1.695 0.495 ;
        RECT  0.360 -0.210 1.525 0.210 ;
        RECT  0.190 -0.210 0.360 0.730 ;
        RECT  0.000 -0.210 0.190 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.725 2.310 1.960 2.730 ;
        RECT  0.555 1.800 0.725 2.730 ;
        RECT  0.000 2.310 0.555 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.635 1.735 1.805 2.165 ;
        RECT  1.085 1.995 1.635 2.115 ;
        RECT  0.915 1.495 1.085 2.115 ;
        RECT  0.360 1.495 0.915 1.615 ;
        RECT  0.190 1.495 0.360 2.075 ;
    END
END AOI22X2AD
MACRO AOI22X4AD
    CLASS CORE ;
    FOREIGN AOI22X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.620 3.290 1.625 ;
        RECT  2.460 0.620 3.150 0.750 ;
        RECT  2.820 1.495 3.150 1.625 ;
        RECT  2.560 1.495 2.820 1.875 ;
        RECT  2.100 1.495 2.560 1.625 ;
        RECT  2.200 0.370 2.460 0.750 ;
        RECT  1.020 0.620 2.200 0.750 ;
        RECT  1.840 1.495 2.100 1.875 ;
        RECT  0.760 0.370 1.020 0.750 ;
        END
        AntennaDiffArea 0.892 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.285 0.870 1.455 1.260 ;
        RECT  0.490 0.870 1.285 0.990 ;
        RECT  0.295 0.870 0.490 1.375 ;
        RECT  0.070 1.145 0.295 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.110 1.160 1.230 ;
        RECT  0.630 1.110 1.050 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.755 0.870 2.900 1.280 ;
        RECT  1.905 0.870 2.755 0.990 ;
        RECT  1.735 0.870 1.905 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 1.110 2.630 1.230 ;
        RECT  2.030 1.110 2.450 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.075 -0.210 3.360 0.210 ;
        RECT  2.905 -0.210 3.075 0.500 ;
        RECT  1.730 -0.210 2.905 0.210 ;
        RECT  1.470 -0.210 1.730 0.500 ;
        RECT  0.365 -0.210 1.470 0.210 ;
        RECT  0.195 -0.210 0.365 0.730 ;
        RECT  0.000 -0.210 0.195 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.335 2.310 3.360 2.730 ;
        RECT  1.165 1.735 1.335 2.730 ;
        RECT  0.615 2.310 1.165 2.730 ;
        RECT  0.445 1.735 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.965 1.745 3.135 2.175 ;
        RECT  2.415 2.020 2.965 2.140 ;
        RECT  2.245 1.745 2.415 2.175 ;
        RECT  1.695 2.020 2.245 2.140 ;
        RECT  1.525 1.495 1.695 2.185 ;
        RECT  0.975 1.495 1.525 1.615 ;
        RECT  0.805 1.495 0.975 2.040 ;
        RECT  0.255 1.495 0.805 1.615 ;
        RECT  0.085 1.495 0.255 2.185 ;
    END
END AOI22X4AD
MACRO AOI22XLAD
    CLASS CORE ;
    FOREIGN AOI22XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.740 1.610 1.660 ;
        RECT  0.895 0.740 1.470 0.860 ;
        RECT  1.040 1.500 1.470 1.660 ;
        RECT  0.725 0.685 0.895 0.860 ;
        END
        AntennaDiffArea 0.162 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.980 0.230 1.435 ;
        END
        AntennaGateArea 0.0604 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.980 0.710 1.375 ;
        END
        AntennaGateArea 0.0603 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.980 1.350 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.845 0.980 1.070 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.535 -0.210 1.680 0.210 ;
        RECT  1.365 -0.210 1.535 0.610 ;
        RECT  0.270 -0.210 1.365 0.210 ;
        RECT  0.100 -0.210 0.270 0.855 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.580 2.310 1.680 2.730 ;
        RECT  0.395 1.530 0.580 2.730 ;
        RECT  0.000 2.310 0.395 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
	 END
END AOI22XLAD
MACRO AOI2B1X1AD
    CLASS CORE ;
    FOREIGN AOI2B1X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.875 0.780 1.890 1.610 ;
        RECT  1.750 0.780 1.875 1.930 ;
        RECT  1.435 0.780 1.750 0.900 ;
        RECT  1.705 1.500 1.750 1.930 ;
        RECT  1.265 0.560 1.435 0.900 ;
        END
        AntennaDiffArea 0.216 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.020 1.630 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.280 1.280 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.0416 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 1.040 1.330 1.375 ;
        END
        AntennaGateArea 0.0904 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.840 -0.210 1.960 0.210 ;
        RECT  1.580 -0.210 1.840 0.660 ;
        RECT  0.815 -0.210 1.580 0.210 ;
        RECT  0.640 -0.210 0.815 0.760 ;
        RECT  0.000 -0.210 0.640 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 2.310 1.960 2.730 ;
        RECT  0.910 2.220 1.170 2.730 ;
        RECT  0.300 2.310 0.910 2.730 ;
        RECT  0.105 1.815 0.300 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.345 1.525 1.515 1.955 ;
        RECT  0.655 1.755 1.345 1.955 ;
        RECT  0.560 1.005 0.950 1.265 ;
        RECT  0.520 1.005 0.560 1.590 ;
        RECT  0.400 0.575 0.520 1.590 ;
        RECT  0.095 0.575 0.400 0.745 ;
    END
END AOI2B1X1AD
MACRO AOI2B1X2AD
    CLASS CORE ;
    FOREIGN AOI2B1X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.070 0.625 2.170 1.690 ;
        RECT  2.030 0.625 2.070 1.975 ;
        RECT  1.660 0.625 2.030 0.745 ;
        RECT  1.900 1.545 2.030 1.975 ;
        RECT  1.400 0.365 1.660 0.745 ;
        END
        AntennaDiffArea 0.41 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.665 0.865 1.890 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.190 1.020 0.380 1.375 ;
        RECT  0.070 1.120 0.190 1.375 ;
        END
        AntennaGateArea 0.0654 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.865 1.480 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.985 -0.210 2.240 0.210 ;
        RECT  1.815 -0.210 1.985 0.495 ;
        RECT  0.875 -0.210 1.815 0.210 ;
        RECT  0.875 0.410 1.035 0.530 ;
        RECT  0.680 -0.210 0.875 0.530 ;
        RECT  0.000 -0.210 0.680 0.210 ;
        RECT  0.515 0.410 0.680 0.530 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.350 2.310 2.240 2.730 ;
        RECT  1.180 1.760 1.350 2.730 ;
        RECT  0.290 2.310 1.180 2.730 ;
        RECT  0.120 1.495 0.290 2.730 ;
        RECT  0.000 2.310 0.120 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.540 1.520 1.710 2.025 ;
        RECT  0.990 1.520 1.540 1.640 ;
        RECT  0.670 1.045 1.070 1.215 ;
        RECT  0.820 1.520 0.990 1.990 ;
        RECT  0.500 0.725 0.670 1.665 ;
        RECT  0.180 0.725 0.500 0.895 ;
    END
END AOI2B1X2AD
MACRO AOI2B1X4AD
    CLASS CORE ;
    FOREIGN AOI2B1X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.200 0.620 3.290 1.550 ;
        RECT  3.150 0.365 3.200 1.550 ;
        RECT  2.940 0.365 3.150 0.745 ;
        RECT  2.795 1.430 3.150 1.550 ;
        RECT  2.370 0.620 2.940 0.745 ;
        RECT  2.625 1.430 2.795 1.885 ;
        RECT  2.110 0.365 2.370 0.745 ;
        RECT  1.090 0.620 2.110 0.745 ;
        RECT  0.830 0.365 1.090 0.745 ;
        END
        AntennaDiffArea 0.754 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.730 1.045 2.915 1.215 ;
        RECT  2.310 0.865 2.730 1.215 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.040 0.375 1.300 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.1298 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.005 0.865 2.150 1.260 ;
        RECT  1.190 0.865 2.005 0.985 ;
        RECT  0.910 0.865 1.190 1.140 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.750 -0.210 3.360 0.210 ;
        RECT  2.580 -0.210 2.750 0.500 ;
        RECT  1.695 -0.210 2.580 0.210 ;
        RECT  1.525 -0.210 1.695 0.500 ;
        RECT  0.305 -0.210 1.525 0.210 ;
        RECT  0.135 -0.210 0.305 0.710 ;
        RECT  0.000 -0.210 0.135 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.075 2.310 3.360 2.730 ;
        RECT  1.905 1.740 2.075 2.730 ;
        RECT  1.355 2.310 1.905 2.730 ;
        RECT  1.185 1.780 1.355 2.730 ;
        RECT  0.255 2.310 1.185 2.730 ;
        RECT  0.085 1.540 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.985 1.710 3.155 2.140 ;
        RECT  2.435 2.020 2.985 2.140 ;
        RECT  2.265 1.500 2.435 2.140 ;
        RECT  1.715 1.500 2.265 1.620 ;
        RECT  1.495 1.140 1.840 1.265 ;
        RECT  1.545 1.500 1.715 2.045 ;
        RECT  0.995 1.500 1.545 1.620 ;
        RECT  1.320 1.140 1.495 1.380 ;
        RECT  0.665 1.260 1.320 1.380 ;
        RECT  0.825 1.500 0.995 1.995 ;
        RECT  0.615 0.460 0.665 1.380 ;
        RECT  0.495 0.460 0.615 1.970 ;
        RECT  0.445 1.540 0.495 1.970 ;
    END
END AOI2B1X4AD
MACRO AOI2B1XLAD
    CLASS CORE ;
    FOREIGN AOI2B1XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.830 1.890 1.815 ;
        RECT  1.435 0.830 1.750 0.950 ;
        RECT  1.705 1.645 1.750 1.815 ;
        RECT  1.265 0.565 1.435 0.950 ;
        END
        AntennaDiffArea 0.144 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.070 1.630 1.470 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.980 0.280 1.240 ;
        RECT  0.070 0.980 0.210 1.655 ;
        END
        AntennaGateArea 0.0404 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.070 1.330 1.470 ;
        END
        AntennaGateArea 0.0604 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.775 -0.210 1.960 0.210 ;
        RECT  1.775 0.590 1.840 0.710 ;
        RECT  1.655 -0.210 1.775 0.710 ;
        RECT  0.810 -0.210 1.655 0.210 ;
        RECT  1.580 0.590 1.655 0.710 ;
        RECT  0.640 -0.210 0.810 0.780 ;
        RECT  0.000 -0.210 0.640 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.135 2.310 1.960 2.730 ;
        RECT  0.965 2.125 1.135 2.730 ;
        RECT  0.300 2.310 0.965 2.730 ;
        RECT  0.105 1.805 0.300 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  0.610 1.710 1.560 1.880 ;
        RECT  0.585 1.055 0.990 1.255 ;
        RECT  0.520 1.055 0.585 1.590 ;
        RECT  0.400 0.565 0.520 1.590 ;
        RECT  0.095 0.565 0.400 0.735 ;
    END
END AOI2B1XLAD
MACRO AOI2BB1X1AD
    CLASS CORE ;
    FOREIGN AOI2BB1X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.540 0.705 1.610 1.655 ;
        RECT  1.490 0.705 1.540 1.945 ;
        RECT  1.060 0.705 1.490 0.825 ;
        RECT  1.420 1.425 1.490 1.945 ;
        END
        AntennaDiffArea 0.241 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 0.980 1.050 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.020 0.770 1.375 ;
        END
        AntennaGateArea 0.0554 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.240 1.300 ;
        END
        AntennaGateArea 0.055 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.565 -0.210 1.680 0.210 ;
        RECT  1.395 -0.210 1.565 0.380 ;
        RECT  0.560 -0.210 1.395 0.210 ;
        RECT  0.560 0.330 0.755 0.450 ;
        RECT  0.440 -0.210 0.560 0.450 ;
        RECT  0.000 -0.210 0.440 0.210 ;
        RECT  0.235 0.330 0.440 0.450 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.915 2.310 1.680 2.730 ;
        RECT  0.745 1.740 0.915 2.730 ;
        RECT  0.000 2.310 0.745 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.290 0.980 1.350 1.265 ;
        RECT  1.170 0.980 1.290 1.615 ;
        RECT  0.480 1.495 1.170 1.615 ;
        RECT  0.480 0.760 0.630 0.880 ;
        RECT  0.360 0.760 0.480 1.615 ;
        RECT  0.255 1.495 0.360 1.615 ;
        RECT  0.085 1.495 0.255 1.665 ;
    END
END AOI2BB1X1AD
MACRO AOI2BB1X2AD
    CLASS CORE ;
    FOREIGN AOI2BB1X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.490 0.675 1.610 2.020 ;
        RECT  1.235 0.675 1.490 0.795 ;
        RECT  1.450 1.425 1.490 2.020 ;
        RECT  1.065 0.365 1.235 0.795 ;
        END
        AntennaDiffArea 0.44 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.915 1.060 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.960 0.790 1.375 ;
        END
        AntennaGateArea 0.073 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.270 1.280 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.0735 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.595 -0.210 1.680 0.210 ;
        RECT  1.425 -0.210 1.595 0.555 ;
        RECT  0.855 -0.210 1.425 0.210 ;
        RECT  0.685 -0.210 0.855 0.415 ;
        RECT  0.255 -0.210 0.685 0.210 ;
        RECT  0.085 -0.210 0.255 0.405 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.935 2.310 1.680 2.730 ;
        RECT  0.765 1.735 0.935 2.730 ;
        RECT  0.000 2.310 0.765 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.300 1.030 1.370 1.290 ;
        RECT  1.180 1.030 1.300 1.615 ;
        RECT  0.510 1.495 1.180 1.615 ;
        RECT  0.510 0.675 0.565 0.845 ;
        RECT  0.390 0.675 0.510 1.615 ;
        RECT  0.255 1.495 0.390 1.615 ;
        RECT  0.085 1.495 0.255 1.670 ;
    END
END AOI2BB1X2AD
MACRO AOI2BB1X4AD
    CLASS CORE ;
    FOREIGN AOI2BB1X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.780 2.450 1.665 ;
        RECT  2.075 0.780 2.310 0.910 ;
        RECT  1.760 1.530 2.310 1.665 ;
        RECT  1.905 0.405 2.075 0.910 ;
        RECT  1.400 0.590 1.905 0.720 ;
        RECT  1.500 1.530 1.760 2.170 ;
        RECT  1.140 0.340 1.400 0.720 ;
        END
        AntennaDiffArea 0.602 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.020 1.030 2.190 1.410 ;
        RECT  1.330 1.290 2.020 1.410 ;
        RECT  1.040 1.090 1.330 1.410 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.090 0.890 1.455 ;
        END
        AntennaGateArea 0.147 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.270 1.280 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.147 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 -0.210 2.520 0.210 ;
        RECT  2.265 -0.210 2.435 0.650 ;
        RECT  1.715 -0.210 2.265 0.210 ;
        RECT  1.545 -0.210 1.715 0.455 ;
        RECT  0.995 -0.210 1.545 0.210 ;
        RECT  0.825 -0.210 0.995 0.700 ;
        RECT  0.275 -0.210 0.825 0.210 ;
        RECT  0.105 -0.210 0.275 0.740 ;
        RECT  0.000 -0.210 0.105 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.325 2.310 2.520 2.730 ;
        RECT  2.155 1.790 2.325 2.730 ;
        RECT  1.045 2.310 2.155 2.730 ;
        RECT  0.875 1.585 1.045 2.730 ;
        RECT  0.000 2.310 0.875 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.450 0.850 1.710 1.170 ;
        RECT  0.635 0.850 1.450 0.970 ;
        RECT  0.510 0.475 0.635 0.970 ;
        RECT  0.465 0.475 0.510 1.765 ;
        RECT  0.390 0.850 0.465 1.765 ;
        RECT  0.375 1.510 0.390 1.765 ;
        RECT  0.205 1.510 0.375 2.070 ;
    END
END AOI2BB1X4AD
MACRO AOI2BB1XLAD
    CLASS CORE ;
    FOREIGN AOI2BB1XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.490 0.735 1.610 1.705 ;
        RECT  1.090 0.735 1.490 0.855 ;
        RECT  1.450 1.425 1.490 1.705 ;
        END
        AntennaDiffArea 0.16 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 1.000 1.070 1.375 ;
        END
        AntennaGateArea 0.0603 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.020 0.770 1.375 ;
        END
        AntennaGateArea 0.0554 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.240 1.300 ;
        END
        AntennaGateArea 0.055 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.565 -0.210 1.680 0.210 ;
        RECT  1.395 -0.210 1.565 0.445 ;
        RECT  0.945 -0.210 1.395 0.210 ;
        RECT  0.775 -0.210 0.945 0.880 ;
        RECT  0.260 -0.210 0.775 0.210 ;
        RECT  0.090 -0.210 0.260 0.445 ;
        RECT  0.000 -0.210 0.090 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.885 2.310 1.680 2.730 ;
        RECT  0.715 1.740 0.885 2.730 ;
        RECT  0.000 2.310 0.715 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.330 1.020 1.370 1.280 ;
        RECT  1.210 1.020 1.330 1.615 ;
        RECT  0.480 1.495 1.210 1.615 ;
        RECT  0.480 0.710 0.585 0.880 ;
        RECT  0.360 0.710 0.480 1.615 ;
        RECT  0.255 1.495 0.360 1.615 ;
        RECT  0.085 1.495 0.255 1.665 ;
    END
END AOI2BB1XLAD
MACRO AOI2BB2X1AD
    CLASS CORE ;
    FOREIGN AOI2BB2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.625 2.170 2.020 ;
        RECT  1.500 0.625 2.030 0.745 ;
        RECT  2.010 1.500 2.030 2.020 ;
        END
        AntennaDiffArea 0.216 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.055 0.865 1.330 1.230 ;
        END
        AntennaGateArea 0.0901 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.865 1.630 1.240 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.230 1.470 ;
        END
        AntennaGateArea 0.0554 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.495 1.025 0.675 1.245 ;
        RECT  0.350 1.025 0.495 1.655 ;
        END
        AntennaGateArea 0.055 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.095 -0.210 2.240 0.210 ;
        RECT  1.925 -0.210 2.095 0.500 ;
        RECT  0.710 -0.210 1.925 0.210 ;
        RECT  0.710 0.330 0.985 0.450 ;
        RECT  0.475 -0.210 0.710 0.450 ;
        RECT  0.000 -0.210 0.475 0.210 ;
        RECT  0.205 0.330 0.475 0.450 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.435 2.310 2.240 2.730 ;
        RECT  1.265 1.850 1.435 2.730 ;
        RECT  0.280 2.310 1.265 2.730 ;
        RECT  0.110 1.955 0.280 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.870 1.040 1.910 1.300 ;
        RECT  1.750 1.040 1.870 1.490 ;
        RECT  1.580 1.610 1.840 1.990 ;
        RECT  0.935 1.370 1.750 1.490 ;
        RECT  1.075 1.610 1.580 1.730 ;
        RECT  0.955 1.610 1.075 2.035 ;
        RECT  0.905 1.865 0.955 2.035 ;
        RECT  0.815 0.735 0.935 1.490 ;
        RECT  0.375 0.735 0.815 0.905 ;
        RECT  0.795 1.370 0.815 1.490 ;
        RECT  0.625 1.370 0.795 1.580 ;
    END
END AOI2BB2X1AD
MACRO AOI2BB2X2AD
    CLASS CORE ;
    FOREIGN AOI2BB2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.155 0.625 2.170 1.740 ;
        RECT  2.030 0.625 2.155 2.055 ;
        RECT  1.760 0.625 2.030 0.745 ;
        RECT  1.985 1.625 2.030 2.055 ;
        RECT  1.500 0.365 1.760 0.745 ;
        END
        AntennaDiffArea 0.394 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.585 1.330 1.250 ;
        RECT  1.055 0.920 1.190 1.250 ;
        END
        AntennaGateArea 0.1629 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.865 1.630 1.250 ;
        END
        AntennaGateArea 0.1629 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.230 1.470 ;
        END
        AntennaGateArea 0.0743 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.495 1.065 0.685 1.245 ;
        RECT  0.350 1.065 0.495 1.655 ;
        END
        AntennaGateArea 0.0745 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.075 -0.210 2.240 0.210 ;
        RECT  1.905 -0.210 2.075 0.495 ;
        RECT  1.020 -0.210 1.905 0.210 ;
        RECT  0.850 -0.210 1.020 0.565 ;
        RECT  0.345 -0.210 0.850 0.210 ;
        RECT  0.175 -0.210 0.345 0.405 ;
        RECT  0.000 -0.210 0.175 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.435 2.310 2.240 2.730 ;
        RECT  1.265 1.850 1.435 2.730 ;
        RECT  0.255 2.310 1.265 2.730 ;
        RECT  0.085 2.065 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.760 1.040 1.900 1.490 ;
        RECT  1.625 1.610 1.795 2.040 ;
        RECT  0.925 1.370 1.760 1.490 ;
        RECT  1.075 1.610 1.625 1.730 ;
        RECT  0.955 1.610 1.075 2.165 ;
        RECT  0.905 1.995 0.955 2.165 ;
        RECT  0.805 0.735 0.925 1.490 ;
        RECT  0.395 0.735 0.805 0.905 ;
        RECT  0.635 1.370 0.805 1.655 ;
    END
END AOI2BB2X2AD
MACRO AOI2BB2X4AD
    CLASS CORE ;
    FOREIGN AOI2BB2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.480 0.365 2.740 0.745 ;
        RECT  2.300 0.625 2.480 0.745 ;
        RECT  2.180 0.625 2.300 0.920 ;
        RECT  1.890 0.800 2.180 0.920 ;
        RECT  1.750 0.800 1.890 1.515 ;
        RECT  1.675 0.800 1.750 0.920 ;
        RECT  1.605 1.395 1.750 1.515 ;
        RECT  1.505 0.390 1.675 0.920 ;
        RECT  1.435 1.395 1.605 1.890 ;
        END
        AntennaDiffArea 0.608 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.025 1.015 3.195 1.410 ;
        RECT  2.205 1.290 3.025 1.410 ;
        RECT  2.030 1.075 2.205 1.410 ;
        END
        AntennaGateArea 0.324 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.735 1.050 2.870 1.170 ;
        RECT  2.440 0.865 2.735 1.170 ;
        RECT  2.350 1.050 2.440 1.170 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.040 1.050 1.375 ;
        END
        AntennaGateArea 0.1479 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.270 1.280 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.147 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.315 -0.210 3.640 0.210 ;
        RECT  3.145 -0.210 3.315 0.785 ;
        RECT  2.060 -0.210 3.145 0.210 ;
        RECT  1.890 -0.210 2.060 0.675 ;
        RECT  1.155 -0.210 1.890 0.210 ;
        RECT  1.155 0.505 1.285 0.675 ;
        RECT  0.980 -0.210 1.155 0.675 ;
        RECT  0.265 -0.210 0.980 0.210 ;
        RECT  0.855 0.505 0.980 0.675 ;
        RECT  0.095 -0.210 0.265 0.745 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.050 2.310 3.640 2.730 ;
        RECT  2.880 1.845 3.050 2.730 ;
        RECT  2.325 2.310 2.880 2.730 ;
        RECT  2.155 1.905 2.325 2.730 ;
        RECT  0.875 2.310 2.155 2.730 ;
        RECT  0.705 1.675 0.875 2.730 ;
        RECT  0.000 2.310 0.705 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  3.240 1.550 3.410 2.025 ;
        RECT  2.685 1.550 3.240 1.685 ;
        RECT  2.515 1.550 2.685 2.015 ;
        RECT  1.965 1.640 2.515 1.760 ;
        RECT  1.795 1.640 1.965 2.140 ;
        RECT  1.245 2.020 1.795 2.140 ;
        RECT  1.385 1.065 1.630 1.235 ;
        RECT  1.225 0.800 1.385 1.235 ;
        RECT  1.075 1.585 1.245 2.140 ;
        RECT  0.630 0.800 1.225 0.920 ;
        RECT  0.510 0.425 0.630 0.920 ;
        RECT  0.460 0.425 0.510 1.670 ;
        RECT  0.390 0.800 0.460 1.670 ;
        RECT  0.265 1.550 0.390 1.670 ;
        RECT  0.095 1.550 0.265 2.025 ;
    END
END AOI2BB2X4AD
MACRO AOI2BB2XLAD
    CLASS CORE ;
    FOREIGN AOI2BB2XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.625 2.170 1.935 ;
        RECT  1.500 0.625 2.030 0.745 ;
        RECT  1.985 1.765 2.030 1.935 ;
        END
        AntennaDiffArea 0.144 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.055 0.865 1.330 1.250 ;
        END
        AntennaGateArea 0.0602 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.865 1.660 1.250 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.230 1.470 ;
        END
        AntennaGateArea 0.0554 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.495 1.025 0.675 1.245 ;
        RECT  0.350 1.025 0.495 1.655 ;
        END
        AntennaGateArea 0.0554 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 -0.210 2.240 0.210 ;
        RECT  1.880 -0.210 2.140 0.505 ;
        RECT  0.740 -0.210 1.880 0.210 ;
        RECT  0.740 0.330 0.985 0.450 ;
        RECT  0.470 -0.210 0.740 0.450 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        RECT  0.205 0.330 0.470 0.450 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.435 2.310 2.240 2.730 ;
        RECT  1.265 1.850 1.435 2.730 ;
        RECT  0.280 2.310 1.265 2.730 ;
        RECT  0.110 1.955 0.280 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.780 1.040 1.900 1.490 ;
        RECT  1.625 1.610 1.795 1.945 ;
        RECT  0.935 1.370 1.780 1.490 ;
        RECT  1.075 1.610 1.625 1.730 ;
        RECT  0.955 1.610 1.075 2.035 ;
        RECT  0.905 1.865 0.955 2.035 ;
        RECT  0.815 0.735 0.935 1.490 ;
        RECT  0.375 0.735 0.815 0.905 ;
        RECT  0.795 1.370 0.815 1.490 ;
        RECT  0.625 1.370 0.795 1.580 ;
    END
END AOI2BB2XLAD
MACRO AOI31X1AD
    CLASS CORE ;
    FOREIGN AOI31X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.780 1.610 1.945 ;
        RECT  1.205 0.780 1.470 0.900 ;
        RECT  1.450 1.425 1.470 1.945 ;
        RECT  1.035 0.710 1.205 0.900 ;
        END
        AntennaDiffArea 0.216 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.020 1.350 1.280 ;
        RECT  1.170 1.020 1.330 1.410 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.030 0.230 1.655 ;
        END
        AntennaGateArea 0.0884 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.980 0.730 1.405 ;
        END
        AntennaGateArea 0.0884 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 1.020 1.050 1.410 ;
        END
        AntennaGateArea 0.0904 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.585 -0.210 1.680 0.210 ;
        RECT  1.415 -0.210 1.585 0.655 ;
        RECT  0.305 -0.210 1.415 0.210 ;
        RECT  0.135 -0.210 0.305 0.860 ;
        RECT  0.000 -0.210 0.135 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.685 2.310 1.680 2.730 ;
        RECT  0.255 2.195 0.685 2.730 ;
        RECT  0.000 2.310 0.255 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.020 1.530 1.280 1.910 ;
        RECT  0.610 1.530 1.020 1.650 ;
        RECT  0.350 1.530 0.610 1.910 ;
    END
END AOI31X1AD
MACRO AOI31X2AD
    CLASS CORE ;
    FOREIGN AOI31X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.780 0.620 1.890 1.590 ;
        RECT  1.730 0.620 1.780 2.115 ;
        RECT  1.360 0.620 1.730 0.740 ;
        RECT  1.585 1.415 1.730 2.115 ;
        RECT  1.100 0.360 1.360 0.740 ;
        END
        AntennaDiffArea 0.394 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.860 1.610 1.260 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.060 0.510 1.230 ;
        RECT  0.070 1.060 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.585 0.865 1.260 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.015 0.865 1.330 1.260 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.675 -0.210 1.960 0.210 ;
        RECT  1.505 -0.210 1.675 0.500 ;
        RECT  0.405 -0.210 1.505 0.210 ;
        RECT  0.235 -0.210 0.405 0.795 ;
        RECT  0.000 -0.210 0.235 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.035 2.310 1.960 2.730 ;
        RECT  0.865 1.695 1.035 2.730 ;
        RECT  0.315 2.310 0.865 2.730 ;
        RECT  0.145 1.525 0.315 2.730 ;
        RECT  0.000 2.310 0.145 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.225 1.405 1.395 2.095 ;
        RECT  0.675 1.405 1.225 1.525 ;
        RECT  0.505 1.405 0.675 2.100 ;
    END
END AOI31X2AD
MACRO AOI31X4AD
    CLASS CORE ;
    FOREIGN AOI31X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.195 0.770 3.290 1.620 ;
        RECT  3.150 0.375 3.195 1.620 ;
        RECT  3.025 0.375 3.150 0.910 ;
        RECT  2.835 1.470 3.150 1.620 ;
        RECT  2.395 0.770 3.025 0.910 ;
        RECT  2.665 1.470 2.835 1.900 ;
        RECT  2.225 0.365 2.395 0.910 ;
        RECT  0.435 0.620 2.225 0.745 ;
        RECT  0.265 0.360 0.435 0.790 ;
        END
        AntennaDiffArea 0.77 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.470 1.045 2.900 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 1.110 1.550 1.230 ;
        RECT  1.145 1.110 1.375 1.330 ;
        RECT  1.030 1.110 1.145 1.230 ;
        END
        AntennaGateArea 0.324 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.685 0.865 1.905 1.260 ;
        RECT  0.900 0.865 1.685 0.985 ;
        RECT  0.630 0.865 0.900 1.260 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.035 1.040 2.205 1.570 ;
        RECT  0.500 1.450 2.035 1.570 ;
        RECT  0.315 1.035 0.500 1.570 ;
        RECT  0.070 1.145 0.315 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.840 -0.210 3.360 0.210 ;
        RECT  2.580 -0.210 2.840 0.650 ;
        RECT  1.440 -0.210 2.580 0.210 ;
        RECT  1.180 -0.210 1.440 0.500 ;
        RECT  0.000 -0.210 1.180 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.115 2.310 3.360 2.730 ;
        RECT  1.945 1.955 2.115 2.730 ;
        RECT  1.395 2.310 1.945 2.730 ;
        RECT  1.225 1.930 1.395 2.730 ;
        RECT  0.675 2.310 1.225 2.730 ;
        RECT  0.505 1.930 0.675 2.730 ;
        RECT  0.000 2.310 0.505 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.980 1.760 3.240 2.140 ;
        RECT  2.475 2.020 2.980 2.140 ;
        RECT  2.305 1.690 2.475 2.140 ;
        RECT  1.755 1.690 2.305 1.810 ;
        RECT  1.585 1.690 1.755 2.135 ;
        RECT  1.035 1.690 1.585 1.810 ;
        RECT  0.865 1.690 1.035 2.120 ;
        RECT  0.315 1.690 0.865 1.810 ;
        RECT  0.145 1.690 0.315 2.120 ;
    END
END AOI31X4AD
MACRO AOI31XLAD
    CLASS CORE ;
    FOREIGN AOI31XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.730 1.610 1.715 ;
        RECT  1.035 0.730 1.470 0.900 ;
        RECT  1.425 1.545 1.470 1.715 ;
        END
        AntennaDiffArea 0.144 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.020 1.350 1.410 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.020 0.230 1.655 ;
        END
        AntennaGateArea 0.0604 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.020 0.730 1.405 ;
        END
        AntennaGateArea 0.0604 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 1.020 1.050 1.410 ;
        END
        AntennaGateArea 0.0604 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.585 -0.210 1.680 0.210 ;
        RECT  1.415 -0.210 1.585 0.610 ;
        RECT  0.305 -0.210 1.415 0.210 ;
        RECT  0.135 -0.210 0.305 0.900 ;
        RECT  0.000 -0.210 0.135 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.590 2.310 1.680 2.730 ;
        RECT  0.590 2.005 0.845 2.175 ;
        RECT  0.390 2.005 0.590 2.730 ;
        RECT  0.155 2.005 0.390 2.175 ;
        RECT  0.000 2.310 0.390 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  0.395 1.530 1.235 1.700 ;
    END
END AOI31XLAD
MACRO AOI32X1AD
    CLASS CORE ;
    FOREIGN AOI32X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.705 2.170 1.640 ;
        RECT  1.300 0.705 2.030 0.825 ;
        RECT  1.775 1.520 2.030 1.640 ;
        RECT  1.515 1.520 1.775 1.900 ;
        RECT  1.130 0.655 1.300 0.825 ;
        END
        AntennaDiffArea 0.27 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.620 0.945 1.890 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.945 1.495 1.375 ;
        END
        AntennaGateArea 0.0906 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.295 1.020 0.470 1.375 ;
        RECT  0.070 1.120 0.295 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.585 0.780 1.300 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.900 0.950 1.070 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.000 -0.210 2.240 0.210 ;
        RECT  1.830 -0.210 2.000 0.585 ;
        RECT  0.320 -0.210 1.830 0.210 ;
        RECT  0.150 -0.210 0.320 0.850 ;
        RECT  0.000 -0.210 0.150 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.010 2.310 2.240 2.730 ;
        RECT  0.815 1.735 1.010 2.730 ;
        RECT  0.285 2.310 0.815 2.730 ;
        RECT  0.115 1.515 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.920 1.775 2.090 2.140 ;
        RECT  1.370 2.020 1.920 2.140 ;
        RECT  1.200 1.495 1.370 2.140 ;
        RECT  0.645 1.495 1.200 1.615 ;
        RECT  0.475 1.495 0.645 1.955 ;
    END
END AOI32X1AD
MACRO AOI32X2AD
    CLASS CORE ;
    FOREIGN AOI32X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.625 2.170 1.640 ;
        RECT  1.360 0.625 2.030 0.745 ;
        RECT  1.740 1.520 2.030 1.640 ;
        RECT  1.480 1.520 1.740 1.900 ;
        RECT  1.100 0.365 1.360 0.745 ;
        END
        AntennaDiffArea 0.504 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.620 0.865 1.890 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.865 1.460 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.030 0.440 1.375 ;
        RECT  0.070 1.145 0.320 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 0.585 0.770 1.280 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 0.865 1.070 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.945 -0.210 2.240 0.210 ;
        RECT  1.775 -0.210 1.945 0.505 ;
        RECT  0.315 -0.210 1.775 0.210 ;
        RECT  0.145 -0.210 0.315 0.840 ;
        RECT  0.000 -0.210 0.145 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.975 2.310 2.240 2.730 ;
        RECT  0.805 1.755 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.500 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.885 1.805 2.055 2.140 ;
        RECT  1.335 2.020 1.885 2.140 ;
        RECT  1.165 1.495 1.335 2.140 ;
        RECT  0.615 1.495 1.165 1.615 ;
        RECT  0.445 1.495 0.615 2.015 ;
    END
END AOI32X2AD
MACRO AOI32X4AD
    CLASS CORE ;
    FOREIGN AOI32X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.990 0.620 4.130 1.680 ;
        RECT  3.300 0.620 3.990 0.790 ;
        RECT  3.690 1.510 3.990 1.680 ;
        RECT  3.430 1.510 3.690 1.890 ;
        RECT  2.970 1.510 3.430 1.680 ;
        RECT  3.130 0.360 3.300 0.790 ;
        RECT  2.090 0.620 3.130 0.790 ;
        RECT  2.710 1.510 2.970 1.890 ;
        RECT  1.920 0.380 2.090 0.790 ;
        RECT  1.205 0.380 1.920 0.550 ;
        END
        AntennaDiffArea 1.01 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.615 1.015 3.790 1.380 ;
        RECT  2.780 1.260 3.615 1.380 ;
        RECT  2.545 0.910 2.780 1.380 ;
        END
        AntennaGateArea 0.324 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.425 1.020 3.470 1.140 ;
        RECT  3.055 0.910 3.425 1.140 ;
        RECT  2.950 1.020 3.055 1.140 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.105 1.000 2.275 1.500 ;
        RECT  0.510 1.380 2.105 1.500 ;
        RECT  0.390 1.020 0.510 1.500 ;
        RECT  0.350 1.145 0.390 1.500 ;
        RECT  0.070 1.145 0.350 1.380 ;
        END
        AntennaGateArea 0.324 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 0.995 1.960 1.260 ;
        RECT  1.680 0.670 1.800 1.260 ;
        RECT  0.870 0.670 1.680 0.790 ;
        RECT  0.770 0.670 0.870 1.260 ;
        RECT  0.630 0.460 0.770 1.260 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.910 1.560 1.155 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.915 -0.210 4.200 0.210 ;
        RECT  3.745 -0.210 3.915 0.455 ;
        RECT  2.560 -0.210 3.745 0.210 ;
        RECT  2.560 0.380 2.730 0.500 ;
        RECT  2.350 -0.210 2.560 0.500 ;
        RECT  0.445 -0.210 2.350 0.210 ;
        RECT  2.210 0.380 2.350 0.500 ;
        RECT  0.275 -0.210 0.445 0.825 ;
        RECT  0.000 -0.210 0.275 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.185 2.310 4.200 2.730 ;
        RECT  2.015 1.865 2.185 2.730 ;
        RECT  1.465 2.310 2.015 2.730 ;
        RECT  1.295 1.870 1.465 2.730 ;
        RECT  0.745 2.310 1.295 2.730 ;
        RECT  0.575 1.865 0.745 2.730 ;
        RECT  0.000 2.310 0.575 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  3.855 1.825 4.025 2.140 ;
        RECT  3.285 2.020 3.855 2.140 ;
        RECT  3.115 1.860 3.285 2.140 ;
        RECT  2.545 2.020 3.115 2.140 ;
        RECT  2.375 1.620 2.545 2.140 ;
        RECT  1.825 1.620 2.375 1.740 ;
        RECT  1.655 1.620 1.825 2.050 ;
        RECT  1.105 1.620 1.655 1.740 ;
        RECT  0.935 1.620 1.105 2.050 ;
        RECT  0.385 1.620 0.935 1.740 ;
        RECT  0.215 1.620 0.385 2.050 ;
    END
END AOI32X4AD
MACRO AOI32XLAD
    CLASS CORE ;
    FOREIGN AOI32XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.770 0.780 1.890 1.935 ;
        RECT  1.200 0.780 1.770 0.900 ;
        RECT  1.735 1.425 1.770 1.935 ;
        RECT  1.415 1.540 1.735 1.710 ;
        RECT  1.080 0.640 1.200 0.900 ;
        END
        AntennaDiffArea 0.162 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.615 1.020 1.650 1.280 ;
        RECT  1.470 1.020 1.615 1.420 ;
        END
        AntennaGateArea 0.0604 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.020 1.350 1.420 ;
        END
        AntennaGateArea 0.0604 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.010 0.230 1.655 ;
        END
        AntennaGateArea 0.0608 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.010 0.720 1.270 ;
        RECT  0.350 1.010 0.490 1.655 ;
        END
        AntennaGateArea 0.0604 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.960 1.020 1.020 1.280 ;
        RECT  0.840 0.585 0.960 1.280 ;
        RECT  0.630 0.585 0.840 0.815 ;
        END
        AntennaGateArea 0.0604 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.855 -0.210 1.960 0.210 ;
        RECT  1.685 -0.210 1.855 0.660 ;
        RECT  0.295 -0.210 1.685 0.210 ;
        RECT  0.125 -0.210 0.295 0.855 ;
        RECT  0.000 -0.210 0.125 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.915 2.310 1.960 2.730 ;
        RECT  0.745 1.510 0.915 2.730 ;
        RECT  0.230 2.310 0.745 2.730 ;
        RECT  0.110 1.970 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
	 END
END AOI32XLAD
MACRO AOI33X1AD
    CLASS CORE ;
    FOREIGN AOI33X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.625 2.450 1.615 ;
        RECT  2.310 0.625 2.415 1.940 ;
        RECT  1.055 0.625 2.310 0.745 ;
        RECT  2.245 1.495 2.310 1.940 ;
        RECT  1.740 1.495 2.245 1.615 ;
        RECT  1.480 1.495 1.740 1.875 ;
        END
        AntennaDiffArea 0.408 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.315 1.015 0.490 1.375 ;
        RECT  0.070 1.135 0.315 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 0.865 0.770 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.865 2.170 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.865 1.890 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.865 1.460 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.315 -0.210 2.520 0.210 ;
        RECT  2.120 -0.210 2.315 0.505 ;
        RECT  0.315 -0.210 2.120 0.210 ;
        RECT  0.145 -0.210 0.315 0.795 ;
        RECT  0.000 -0.210 0.145 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.000 2.310 2.520 2.730 ;
        RECT  0.780 1.750 1.000 2.730 ;
        RECT  0.255 2.310 0.780 2.730 ;
        RECT  0.085 1.585 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.885 1.770 2.055 2.130 ;
        RECT  1.335 2.010 1.885 2.130 ;
        RECT  1.165 1.495 1.335 2.130 ;
        RECT  0.615 1.495 1.165 1.615 ;
        RECT  0.445 1.495 0.615 1.945 ;
    END
END AOI33X1AD
MACRO AOI33X2AD
    CLASS CORE ;
    FOREIGN AOI33X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.625 2.450 1.615 ;
        RECT  2.310 0.625 2.415 2.185 ;
        RECT  1.335 0.625 2.310 0.745 ;
        RECT  2.245 1.495 2.310 2.185 ;
        RECT  1.740 1.495 2.245 1.615 ;
        RECT  1.480 1.495 1.740 1.875 ;
        RECT  1.075 0.365 1.335 0.745 ;
        END
        AntennaDiffArea 0.76 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 1.020 0.490 1.375 ;
        RECT  0.070 1.115 0.310 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.615 0.760 0.770 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.895 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.865 2.170 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 0.865 1.890 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.865 1.520 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.300 -0.210 2.520 0.210 ;
        RECT  2.100 -0.210 2.300 0.500 ;
        RECT  0.315 -0.210 2.100 0.210 ;
        RECT  0.145 -0.210 0.315 0.795 ;
        RECT  0.000 -0.210 0.145 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.975 2.310 2.520 2.730 ;
        RECT  0.805 1.750 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.615 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.885 1.740 2.055 2.170 ;
        RECT  1.335 2.020 1.885 2.140 ;
        RECT  1.165 1.495 1.335 2.140 ;
        RECT  0.615 1.495 1.165 1.615 ;
        RECT  0.445 1.495 0.615 1.960 ;
    END
END AOI33X2AD
MACRO AOI33X4AD
    CLASS CORE ;
    FOREIGN AOI33X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 0.770 4.690 1.815 ;
        RECT  4.140 0.770 4.530 0.900 ;
        RECT  2.605 1.645 4.530 1.815 ;
        RECT  3.980 0.380 4.140 0.900 ;
        RECT  2.660 0.380 3.980 0.550 ;
        RECT  2.530 0.380 2.660 0.745 ;
        RECT  1.920 0.620 2.530 0.745 ;
        RECT  1.790 0.380 1.920 0.745 ;
        RECT  1.130 0.380 1.790 0.550 ;
        END
        AntennaDiffArea 1.32 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.040 2.160 1.500 ;
        RECT  0.490 1.380 2.000 1.500 ;
        RECT  0.315 1.020 0.490 1.500 ;
        RECT  0.290 1.020 0.315 1.375 ;
        RECT  0.070 1.130 0.290 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.665 1.000 1.820 1.260 ;
        RECT  1.540 0.670 1.665 1.260 ;
        RECT  0.770 0.670 1.540 0.790 ;
        RECT  0.620 0.580 0.770 1.260 ;
        END
        AntennaGateArea 0.324 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.900 0.910 1.420 1.170 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.165 1.020 4.335 1.500 ;
        RECT  2.540 1.380 4.165 1.500 ;
        RECT  2.310 0.865 2.540 1.500 ;
        END
        AntennaGateArea 0.324 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.855 1.095 4.040 1.215 ;
        RECT  3.735 0.670 3.855 1.215 ;
        RECT  3.010 0.670 3.735 0.790 ;
        RECT  2.780 0.670 3.010 1.260 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.135 0.910 3.615 1.195 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.500 -0.210 4.760 0.210 ;
        RECT  4.260 -0.210 4.500 0.555 ;
        RECT  2.390 -0.210 4.260 0.210 ;
        RECT  2.215 -0.210 2.390 0.500 ;
        RECT  0.315 -0.210 2.215 0.210 ;
        RECT  0.145 -0.210 0.315 0.835 ;
        RECT  0.000 -0.210 0.145 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.100 2.310 4.760 2.730 ;
        RECT  1.840 1.870 2.100 2.730 ;
        RECT  1.380 2.310 1.840 2.730 ;
        RECT  1.120 1.870 1.380 2.730 ;
        RECT  0.660 2.310 1.120 2.730 ;
        RECT  0.400 1.870 0.660 2.730 ;
        RECT  0.000 2.310 0.400 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.760 2.520 ;
        LAYER M1 ;
        RECT  4.405 1.955 4.575 2.140 ;
        RECT  3.855 2.020 4.405 2.140 ;
        RECT  3.685 1.970 3.855 2.140 ;
        RECT  3.135 2.020 3.685 2.140 ;
        RECT  2.965 1.970 3.135 2.140 ;
        RECT  2.415 2.020 2.965 2.140 ;
        RECT  2.245 1.620 2.415 2.140 ;
        RECT  1.695 1.620 2.245 1.740 ;
        RECT  1.525 1.620 1.695 2.050 ;
        RECT  0.975 1.620 1.525 1.740 ;
        RECT  0.805 1.620 0.975 2.050 ;
        RECT  0.255 1.620 0.805 1.740 ;
        RECT  0.085 1.620 0.255 2.065 ;
    END
END AOI33X4AD
MACRO AOI33XLAD
    CLASS CORE ;
    FOREIGN AOI33XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.625 2.450 1.630 ;
        RECT  2.310 0.625 2.415 1.790 ;
        RECT  1.055 0.625 2.310 0.745 ;
        RECT  2.245 1.510 2.310 1.790 ;
        RECT  1.695 1.510 2.245 1.630 ;
        RECT  1.515 1.510 1.695 1.825 ;
        END
        AntennaDiffArea 0.272 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.130 0.490 1.390 ;
        RECT  0.320 0.870 0.440 1.390 ;
        RECT  0.070 1.130 0.320 1.390 ;
        END
        AntennaGateArea 0.06 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 0.865 0.770 1.390 ;
        END
        AntennaGateArea 0.06 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.865 1.050 1.390 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.865 2.170 1.390 ;
        END
        AntennaGateArea 0.06 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.810 0.865 1.890 1.115 ;
        RECT  1.650 0.865 1.810 1.390 ;
        END
        AntennaGateArea 0.06 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 0.865 1.460 1.390 ;
        RECT  1.190 1.115 1.320 1.390 ;
        END
        AntennaGateArea 0.06 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.325 -0.210 2.520 0.210 ;
        RECT  2.155 -0.210 2.325 0.500 ;
        RECT  0.315 -0.210 2.155 0.210 ;
        RECT  0.315 0.625 0.360 0.745 ;
        RECT  0.145 -0.210 0.315 0.745 ;
        RECT  0.000 -0.210 0.145 0.210 ;
        RECT  0.100 0.625 0.145 0.745 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.970 2.310 2.520 2.730 ;
        RECT  0.970 1.750 1.020 1.870 ;
        RECT  0.805 1.750 0.970 2.730 ;
        RECT  0.760 1.750 0.805 1.870 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.615 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.840 1.750 2.100 2.130 ;
        RECT  1.335 2.010 1.840 2.130 ;
        RECT  1.165 1.510 1.335 2.130 ;
        RECT  0.615 1.510 1.165 1.630 ;
        RECT  0.445 1.510 0.615 1.770 ;
    END
END AOI33XLAD
MACRO BENCX1AD
    CLASS CORE ;
    FOREIGN BENCX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.755 0.755 7.890 1.610 ;
        RECT  7.745 0.755 7.755 0.880 ;
        RECT  7.585 1.395 7.755 1.610 ;
        RECT  7.575 0.710 7.745 0.880 ;
        END
        AntennaDiffArea 0.364 ;
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.990 0.765 11.130 1.510 ;
        RECT  10.690 0.765 10.990 0.885 ;
        RECT  10.715 1.385 10.990 1.510 ;
        RECT  10.565 1.385 10.715 1.995 ;
        RECT  10.570 0.330 10.690 0.885 ;
        RECT  10.540 1.565 10.565 1.995 ;
        END
        AntennaDiffArea 0.364 ;
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.425 1.750 8.720 2.090 ;
        RECT  5.690 1.970 8.425 2.090 ;
        RECT  5.570 1.835 5.690 2.090 ;
        RECT  4.760 1.835 5.570 1.955 ;
        RECT  4.640 1.835 4.760 2.090 ;
        RECT  3.535 1.970 4.640 2.090 ;
        END
        AntennaGateArea 0.0911 ;
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.185 1.630 4.355 1.845 ;
        RECT  3.325 1.630 4.185 1.750 ;
        RECT  3.205 1.535 3.325 1.750 ;
        RECT  2.450 1.535 3.205 1.655 ;
        RECT  2.310 1.240 2.450 1.655 ;
        RECT  2.105 1.240 2.310 1.360 ;
        END
        AntennaGateArea 0.161 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.470 0.380 4.590 1.110 ;
        RECT  3.335 0.380 4.470 0.500 ;
        RECT  3.215 0.380 3.335 1.120 ;
        RECT  1.955 1.000 3.215 1.120 ;
        RECT  1.835 1.000 1.955 1.375 ;
        RECT  1.750 1.145 1.835 1.375 ;
        END
        AntennaGateArea 0.1464 ;
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.460 1.350 0.680 2.030 ;
        RECT  0.540 0.395 0.660 0.915 ;
        RECT  0.250 0.795 0.540 0.915 ;
        RECT  0.250 1.350 0.460 1.470 ;
        RECT  0.130 0.795 0.250 1.470 ;
        RECT  0.070 1.145 0.130 1.375 ;
        END
        AntennaDiffArea 0.392 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.075 -0.210 11.200 0.210 ;
        RECT  10.905 -0.210 11.075 0.630 ;
        RECT  10.380 -0.210 10.905 0.210 ;
        RECT  10.120 -0.210 10.380 0.300 ;
        RECT  9.855 -0.210 10.120 0.210 ;
        RECT  9.595 -0.210 9.855 0.300 ;
        RECT  9.075 -0.210 9.595 0.210 ;
        RECT  8.815 -0.210 9.075 0.330 ;
        RECT  8.170 -0.210 8.815 0.210 ;
        RECT  7.910 -0.210 8.170 0.310 ;
        RECT  7.410 -0.210 7.910 0.210 ;
        RECT  7.150 -0.210 7.410 0.310 ;
        RECT  5.310 -0.210 7.150 0.210 ;
        RECT  5.050 -0.210 5.310 0.310 ;
        RECT  4.015 -0.210 5.050 0.210 ;
        RECT  3.755 -0.210 4.015 0.260 ;
        RECT  2.505 -0.210 3.755 0.210 ;
        RECT  2.245 -0.210 2.505 0.310 ;
        RECT  1.745 -0.210 2.245 0.210 ;
        RECT  1.485 -0.210 1.745 0.310 ;
        RECT  1.100 -0.210 1.485 0.210 ;
        RECT  0.840 -0.210 1.100 0.510 ;
        RECT  0.320 -0.210 0.840 0.210 ;
        RECT  0.160 -0.210 0.320 0.665 ;
        RECT  0.000 -0.210 0.160 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.065 2.310 11.200 2.730 ;
        RECT  10.915 1.635 11.065 2.730 ;
        RECT  10.380 2.310 10.915 2.730 ;
        RECT  10.120 2.210 10.380 2.730 ;
        RECT  9.105 2.310 10.120 2.730 ;
        RECT  8.845 1.710 9.105 2.730 ;
        RECT  8.315 2.310 8.845 2.730 ;
        RECT  8.055 2.210 8.315 2.730 ;
        RECT  7.555 2.310 8.055 2.730 ;
        RECT  7.295 2.210 7.555 2.730 ;
        RECT  5.320 2.310 7.295 2.730 ;
        RECT  5.060 2.075 5.320 2.730 ;
        RECT  4.100 2.310 5.060 2.730 ;
        RECT  3.840 2.210 4.100 2.730 ;
        RECT  2.580 2.310 3.840 2.730 ;
        RECT  2.060 2.210 2.580 2.730 ;
        RECT  1.100 2.310 2.060 2.730 ;
        RECT  0.840 2.020 1.100 2.730 ;
        RECT  0.290 2.310 0.840 2.730 ;
        RECT  0.170 1.600 0.290 2.730 ;
        RECT  0.000 2.310 0.170 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.200 2.520 ;
        LAYER M1 ;
        RECT  10.445 1.005 10.800 1.265 ;
        RECT  10.325 0.785 10.445 1.480 ;
        RECT  10.020 0.785 10.325 0.905 ;
        RECT  10.020 1.350 10.325 1.480 ;
        RECT  9.760 1.045 10.205 1.215 ;
        RECT  9.900 0.645 10.020 0.905 ;
        RECT  9.900 1.350 10.020 1.870 ;
        RECT  9.695 0.735 9.760 1.580 ;
        RECT  9.640 0.735 9.695 1.655 ;
        RECT  8.570 0.735 9.640 0.855 ;
        RECT  9.525 1.460 9.640 1.655 ;
        RECT  8.715 1.460 9.525 1.580 ;
        RECT  9.400 0.975 9.520 1.340 ;
        RECT  8.140 0.975 9.400 1.095 ;
        RECT  9.275 0.355 9.395 0.615 ;
        RECT  8.380 0.495 9.275 0.615 ;
        RECT  8.305 1.215 9.245 1.335 ;
        RECT  8.455 1.460 8.715 1.630 ;
        RECT  8.260 0.495 8.380 0.855 ;
        RECT  8.185 1.215 8.305 1.850 ;
        RECT  6.205 1.730 8.185 1.850 ;
        RECT  8.020 0.430 8.140 1.095 ;
        RECT  6.720 0.430 8.020 0.550 ;
        RECT  7.125 1.000 7.635 1.260 ;
        RECT  7.005 0.670 7.125 1.590 ;
        RECT  6.840 0.670 7.005 0.930 ;
        RECT  6.720 1.395 6.835 1.600 ;
        RECT  6.600 0.430 6.720 1.600 ;
        RECT  6.465 0.430 6.600 0.550 ;
        RECT  6.575 1.395 6.600 1.600 ;
        RECT  6.455 0.880 6.480 1.140 ;
        RECT  6.205 0.430 6.465 0.760 ;
        RECT  6.335 0.880 6.455 1.465 ;
        RECT  6.080 0.880 6.335 1.000 ;
        RECT  6.230 1.295 6.335 1.465 ;
        RECT  5.315 0.430 6.205 0.550 ;
        RECT  6.065 1.690 6.205 1.850 ;
        RECT  5.700 1.320 6.085 1.440 ;
        RECT  5.960 0.670 6.080 1.000 ;
        RECT  5.945 1.595 6.065 1.850 ;
        RECT  5.820 0.670 5.960 0.790 ;
        RECT  4.595 1.595 5.945 1.715 ;
        RECT  5.580 0.670 5.700 1.440 ;
        RECT  5.435 0.670 5.580 0.790 ;
        RECT  5.405 1.320 5.580 1.440 ;
        RECT  5.315 0.910 5.410 1.170 ;
        RECT  5.195 0.430 5.315 1.170 ;
        RECT  4.885 1.050 5.195 1.170 ;
        RECT  4.860 1.050 4.885 1.460 ;
        RECT  4.740 0.570 4.860 1.460 ;
        RECT  4.715 1.290 4.740 1.460 ;
        RECT  4.475 1.325 4.595 1.715 ;
        RECT  4.350 1.325 4.475 1.445 ;
        RECT  4.230 0.635 4.350 1.445 ;
        RECT  4.180 0.635 4.230 0.805 ;
        RECT  3.580 1.240 3.640 1.470 ;
        RECT  3.580 0.635 3.630 0.805 ;
        RECT  3.460 0.635 3.580 1.470 ;
        RECT  2.575 1.240 3.460 1.360 ;
        RECT  3.020 0.695 3.070 0.865 ;
        RECT  2.900 0.500 3.020 0.865 ;
        RECT  1.830 1.855 2.960 1.975 ;
        RECT  2.125 0.500 2.900 0.620 ;
        RECT  1.710 0.740 2.755 0.860 ;
        RECT  1.865 0.430 2.125 0.620 ;
        RECT  1.660 1.535 1.830 1.975 ;
        RECT  1.590 0.740 1.710 0.995 ;
        RECT  1.380 1.535 1.660 1.655 ;
        RECT  1.380 0.875 1.590 0.995 ;
        RECT  1.265 0.585 1.435 0.755 ;
        RECT  1.290 1.780 1.410 2.080 ;
        RECT  1.260 0.875 1.380 1.655 ;
        RECT  0.990 1.780 1.290 1.900 ;
        RECT  0.990 0.630 1.265 0.755 ;
        RECT  1.140 1.005 1.260 1.525 ;
        RECT  0.870 0.630 0.990 1.900 ;
        RECT  0.375 1.045 0.870 1.215 ;
    END
END BENCX1AD
MACRO BENCX2AD
    CLASS CORE ;
    FOREIGN BENCX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.735 1.400 9.890 1.520 ;
        RECT  9.735 0.750 9.850 0.870 ;
        RECT  9.590 0.750 9.735 1.520 ;
        RECT  8.870 0.750 9.590 0.870 ;
        RECT  8.870 1.400 9.590 1.520 ;
        END
        AntennaDiffArea 0.844 ;
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.385 0.385 13.555 2.105 ;
        RECT  13.370 0.705 13.385 2.105 ;
        RECT  13.230 0.705 13.370 1.535 ;
        RECT  12.855 0.705 13.230 0.880 ;
        RECT  12.860 1.375 13.230 1.535 ;
        RECT  12.690 1.375 12.860 2.105 ;
        RECT  12.690 0.340 12.855 0.880 ;
        END
        AntennaDiffArea 0.844 ;
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.570 1.500 10.775 1.620 ;
        RECT  10.420 1.500 10.570 2.000 ;
        RECT  8.305 1.880 10.420 2.000 ;
        RECT  8.185 1.880 8.305 2.105 ;
        RECT  5.790 1.985 8.185 2.105 ;
        RECT  5.655 1.960 5.790 2.105 ;
        RECT  4.170 1.960 5.655 2.080 ;
        END
        AntennaGateArea 0.1322 ;
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.855 1.670 6.025 1.840 ;
        RECT  3.290 1.720 5.855 1.840 ;
        RECT  3.150 1.215 3.290 1.840 ;
        RECT  3.030 1.215 3.150 1.335 ;
        END
        AntennaGateArea 0.3087 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.770 0.975 4.940 1.145 ;
        RECT  4.570 0.975 4.770 1.095 ;
        RECT  4.450 0.380 4.570 1.095 ;
        RECT  4.075 0.380 4.450 0.500 ;
        RECT  3.955 0.380 4.075 1.095 ;
        RECT  3.665 0.910 3.955 1.095 ;
        RECT  2.680 0.975 3.665 1.095 ;
        RECT  2.560 0.975 2.680 1.270 ;
        RECT  2.510 1.100 2.560 1.270 ;
        END
        AntennaGateArea 0.3098 ;
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 0.340 1.340 0.910 ;
        RECT  1.140 1.360 1.310 2.050 ;
        RECT  0.640 1.360 1.140 1.500 ;
        RECT  0.590 0.790 1.120 0.910 ;
        RECT  0.545 1.360 0.640 2.050 ;
        RECT  0.545 0.340 0.590 0.910 ;
        RECT  0.425 0.340 0.545 2.050 ;
        RECT  0.420 0.340 0.425 1.375 ;
        RECT  0.350 1.145 0.420 1.375 ;
        END
        AntennaDiffArea 0.844 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.890 -0.210 14.000 0.210 ;
        RECT  13.720 -0.210 13.890 0.860 ;
        RECT  13.195 -0.210 13.720 0.210 ;
        RECT  13.025 -0.210 13.195 0.560 ;
        RECT  12.520 -0.210 13.025 0.210 ;
        RECT  12.260 -0.210 12.520 0.680 ;
        RECT  11.755 -0.210 12.260 0.210 ;
        RECT  11.555 -0.210 11.755 0.590 ;
        RECT  10.210 -0.210 11.555 0.210 ;
        RECT  9.950 -0.210 10.210 0.390 ;
        RECT  9.490 -0.210 9.950 0.210 ;
        RECT  9.230 -0.210 9.490 0.390 ;
        RECT  8.770 -0.210 9.230 0.210 ;
        RECT  8.510 -0.210 8.770 0.390 ;
        RECT  7.970 -0.210 8.510 0.210 ;
        RECT  7.710 -0.210 7.970 0.390 ;
        RECT  5.620 -0.210 7.710 0.210 ;
        RECT  5.360 -0.210 5.620 0.300 ;
        RECT  4.865 -0.210 5.360 0.210 ;
        RECT  4.690 -0.210 4.865 0.785 ;
        RECT  3.225 -0.210 4.690 0.210 ;
        RECT  2.965 -0.210 3.225 0.370 ;
        RECT  2.455 -0.210 2.965 0.210 ;
        RECT  2.270 -0.210 2.455 0.545 ;
        RECT  1.740 -0.210 2.270 0.210 ;
        RECT  1.480 -0.210 1.740 0.680 ;
        RECT  1.000 -0.210 1.480 0.210 ;
        RECT  0.780 -0.210 1.000 0.665 ;
        RECT  0.230 -0.210 0.780 0.210 ;
        RECT  0.110 -0.210 0.230 0.860 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.890 2.310 14.000 2.730 ;
        RECT  13.730 1.585 13.890 2.730 ;
        RECT  13.195 2.310 13.730 2.730 ;
        RECT  13.025 1.660 13.195 2.730 ;
        RECT  12.480 2.310 13.025 2.730 ;
        RECT  12.310 1.690 12.480 2.730 ;
        RECT  11.720 2.310 12.310 2.730 ;
        RECT  11.550 1.705 11.720 2.730 ;
        RECT  10.580 2.310 11.550 2.730 ;
        RECT  10.060 2.130 10.580 2.730 ;
        RECT  9.510 2.310 10.060 2.730 ;
        RECT  9.250 2.130 9.510 2.730 ;
        RECT  8.770 2.310 9.250 2.730 ;
        RECT  8.510 2.130 8.770 2.730 ;
        RECT  7.970 2.310 8.510 2.730 ;
        RECT  7.710 2.225 7.970 2.730 ;
        RECT  5.490 2.310 7.710 2.730 ;
        RECT  5.230 2.200 5.490 2.730 ;
        RECT  4.725 2.310 5.230 2.730 ;
        RECT  4.465 2.200 4.725 2.730 ;
        RECT  3.470 2.310 4.465 2.730 ;
        RECT  3.210 2.220 3.470 2.730 ;
        RECT  2.390 2.310 3.210 2.730 ;
        RECT  2.200 1.690 2.390 2.730 ;
        RECT  1.695 2.310 2.200 2.730 ;
        RECT  1.525 1.605 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.800 1.655 0.975 2.730 ;
        RECT  0.255 2.310 0.800 2.730 ;
        RECT  0.085 1.490 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 14.000 2.520 ;
        LAYER M1 ;
        RECT  12.570 1.060 13.095 1.180 ;
        RECT  12.450 0.800 12.570 1.520 ;
        RECT  12.115 0.800 12.450 0.920 ;
        RECT  12.115 1.400 12.450 1.520 ;
        RECT  11.945 0.665 12.115 0.920 ;
        RECT  11.945 1.400 12.115 1.845 ;
        RECT  11.775 1.045 12.100 1.215 ;
        RECT  11.655 0.710 11.775 1.560 ;
        RECT  10.765 0.710 11.655 0.830 ;
        RECT  11.065 1.440 11.655 1.560 ;
        RECT  11.380 0.950 11.500 1.265 ;
        RECT  10.620 0.470 11.420 0.590 ;
        RECT  10.130 0.950 11.380 1.070 ;
        RECT  10.130 1.200 11.230 1.320 ;
        RECT  10.895 1.440 11.065 1.940 ;
        RECT  10.450 0.470 10.620 0.640 ;
        RECT  10.010 0.510 10.130 1.070 ;
        RECT  10.010 1.200 10.130 1.760 ;
        RECT  7.590 0.510 10.010 0.630 ;
        RECT  8.035 1.640 10.010 1.760 ;
        RECT  8.750 1.040 9.405 1.210 ;
        RECT  8.630 0.760 8.750 1.520 ;
        RECT  8.110 0.760 8.630 0.880 ;
        RECT  8.130 1.400 8.630 1.520 ;
        RECT  7.990 1.060 8.510 1.240 ;
        RECT  7.915 1.640 8.035 1.860 ;
        RECT  7.780 1.120 7.990 1.240 ;
        RECT  6.540 1.740 7.915 1.860 ;
        RECT  7.660 1.120 7.780 1.620 ;
        RECT  6.780 1.500 7.660 1.620 ;
        RECT  7.445 0.510 7.590 0.685 ;
        RECT  7.445 1.260 7.515 1.380 ;
        RECT  7.325 0.510 7.445 1.380 ;
        RECT  6.900 0.910 7.325 1.030 ;
        RECT  7.255 1.260 7.325 1.380 ;
        RECT  6.240 0.380 6.980 0.500 ;
        RECT  6.660 0.620 6.780 1.620 ;
        RECT  6.360 0.620 6.660 0.740 ;
        RECT  6.420 0.910 6.540 1.860 ;
        RECT  6.240 0.910 6.420 1.030 ;
        RECT  6.180 1.425 6.300 1.855 ;
        RECT  6.120 0.380 6.240 1.030 ;
        RECT  5.955 1.425 6.180 1.545 ;
        RECT  5.610 0.420 6.120 0.540 ;
        RECT  5.835 0.660 5.955 1.545 ;
        RECT  5.785 0.660 5.835 0.830 ;
        RECT  5.655 1.375 5.835 1.545 ;
        RECT  5.610 1.005 5.705 1.175 ;
        RECT  5.490 0.420 5.610 1.175 ;
        RECT  5.195 1.005 5.490 1.175 ;
        RECT  5.075 0.580 5.195 1.565 ;
        RECT  5.025 0.580 5.075 0.750 ;
        RECT  4.890 1.395 5.075 1.565 ;
        RECT  4.265 0.620 4.330 1.420 ;
        RECT  4.210 0.620 4.265 1.555 ;
        RECT  4.095 1.300 4.210 1.555 ;
        RECT  3.525 1.300 4.095 1.420 ;
        RECT  3.690 1.980 3.860 2.150 ;
        RECT  3.715 0.490 3.835 0.750 ;
        RECT  2.585 0.490 3.715 0.610 ;
        RECT  2.755 1.980 3.690 2.100 ;
        RECT  2.305 0.735 3.545 0.855 ;
        RECT  2.585 1.450 2.755 2.100 ;
        RECT  2.305 1.450 2.585 1.570 ;
        RECT  2.185 0.735 2.305 1.570 ;
        RECT  1.850 1.080 2.185 1.200 ;
        RECT  1.900 1.330 2.045 1.925 ;
        RECT  1.900 0.570 2.030 0.930 ;
        RECT  1.580 0.810 1.900 0.930 ;
        RECT  1.580 1.330 1.900 1.450 ;
        RECT  1.460 0.810 1.580 1.450 ;
        RECT  0.665 1.050 1.460 1.170 ;
    END
END BENCX2AD
MACRO BENCX4AD
    CLASS CORE ;
    FOREIGN BENCX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.625 0.755 14.900 1.520 ;
        RECT  12.360 0.755 14.625 0.875 ;
        RECT  12.360 1.400 14.625 1.520 ;
        END
        AntennaDiffArea 1.688 ;
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  21.180 0.345 21.300 2.055 ;
        RECT  21.025 0.765 21.180 1.535 ;
        RECT  20.580 0.765 21.025 0.925 ;
        RECT  20.580 1.380 21.025 1.535 ;
        RECT  20.460 0.345 20.580 0.925 ;
        RECT  20.460 1.380 20.580 2.055 ;
        RECT  19.885 0.765 20.460 0.925 ;
        RECT  19.905 1.380 20.460 1.535 ;
        RECT  19.740 1.380 19.905 2.065 ;
        RECT  19.860 0.390 19.885 0.925 ;
        RECT  19.740 0.345 19.860 0.925 ;
        RECT  19.715 0.390 19.740 0.925 ;
        RECT  19.230 1.380 19.740 1.535 ;
        RECT  19.140 0.765 19.715 0.925 ;
        RECT  19.020 1.380 19.230 2.055 ;
        RECT  19.020 0.345 19.140 0.925 ;
        END
        AntennaDiffArea 1.688 ;
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  15.495 1.880 15.655 2.170 ;
        RECT  15.425 1.570 15.495 2.170 ;
        RECT  15.325 1.570 15.425 2.000 ;
        RECT  11.855 1.880 15.325 2.000 ;
        RECT  11.735 1.880 11.855 2.100 ;
        RECT  6.455 1.980 11.735 2.100 ;
        END
        AntennaGateArea 0.1934 ;
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.685 1.660 8.855 1.830 ;
        RECT  6.440 1.710 8.685 1.830 ;
        RECT  6.320 1.535 6.440 1.830 ;
        RECT  5.710 1.535 6.320 1.655 ;
        RECT  5.390 1.245 5.710 1.655 ;
        RECT  4.730 1.535 5.390 1.655 ;
        RECT  4.610 1.135 4.730 1.655 ;
        RECT  4.570 1.135 4.610 1.395 ;
        END
        AntennaGateArea 0.5647 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.010 0.520 7.230 1.245 ;
        RECT  6.430 0.520 7.010 0.640 ;
        RECT  6.310 0.520 6.430 1.125 ;
        RECT  5.210 1.005 6.310 1.125 ;
        RECT  5.205 1.005 5.210 1.285 ;
        RECT  5.090 1.005 5.205 1.365 ;
        RECT  4.945 1.245 5.090 1.365 ;
        END
        AntennaGateArea 0.539 ;
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 0.340 2.780 0.910 ;
        RECT  2.580 1.360 2.750 2.050 ;
        RECT  2.030 1.360 2.580 1.515 ;
        RECT  2.080 0.790 2.560 0.910 ;
        RECT  1.860 0.340 2.080 0.910 ;
        RECT  1.850 1.360 2.030 2.050 ;
        RECT  1.310 0.790 1.860 0.910 ;
        RECT  1.310 1.360 1.850 1.515 ;
        RECT  1.190 0.340 1.310 0.910 ;
        RECT  1.190 1.360 1.310 2.000 ;
        RECT  0.690 0.790 1.190 0.910 ;
        RECT  0.690 1.360 1.190 1.515 ;
        RECT  0.590 0.790 0.690 1.515 ;
        RECT  0.470 0.340 0.590 2.020 ;
        RECT  0.380 0.790 0.470 1.515 ;
        RECT  0.350 1.005 0.380 1.515 ;
        END
        AntennaDiffArea 1.688 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  21.680 -0.210 21.840 0.210 ;
        RECT  21.520 -0.210 21.680 0.635 ;
        RECT  20.965 -0.210 21.520 0.210 ;
        RECT  20.795 -0.210 20.965 0.635 ;
        RECT  20.245 -0.210 20.795 0.210 ;
        RECT  20.075 -0.210 20.245 0.635 ;
        RECT  19.525 -0.210 20.075 0.210 ;
        RECT  19.355 -0.210 19.525 0.635 ;
        RECT  18.850 -0.210 19.355 0.210 ;
        RECT  18.590 -0.210 18.850 0.615 ;
        RECT  18.130 -0.210 18.590 0.210 ;
        RECT  17.870 -0.210 18.130 0.585 ;
        RECT  17.160 -0.210 17.870 0.210 ;
        RECT  16.900 -0.210 17.160 0.390 ;
        RECT  16.430 -0.210 16.900 0.210 ;
        RECT  16.170 -0.210 16.430 0.390 ;
        RECT  15.260 -0.210 16.170 0.210 ;
        RECT  15.000 -0.210 15.260 0.390 ;
        RECT  14.520 -0.210 15.000 0.210 ;
        RECT  14.260 -0.210 14.520 0.390 ;
        RECT  13.760 -0.210 14.260 0.210 ;
        RECT  13.500 -0.210 13.760 0.390 ;
        RECT  13.000 -0.210 13.500 0.210 ;
        RECT  12.740 -0.210 13.000 0.390 ;
        RECT  12.240 -0.210 12.740 0.210 ;
        RECT  11.980 -0.210 12.240 0.390 ;
        RECT  11.500 -0.210 11.980 0.210 ;
        RECT  11.240 -0.210 11.500 0.390 ;
        RECT  10.750 -0.210 11.240 0.210 ;
        RECT  10.490 -0.210 10.750 0.745 ;
        RECT  8.050 -0.210 10.490 0.210 ;
        RECT  7.790 -0.210 8.050 0.390 ;
        RECT  7.250 -0.210 7.790 0.210 ;
        RECT  6.990 -0.210 7.250 0.390 ;
        RECT  5.470 -0.210 6.990 0.210 ;
        RECT  5.210 -0.210 5.470 0.400 ;
        RECT  3.900 -0.210 5.210 0.210 ;
        RECT  3.640 -0.210 3.900 0.590 ;
        RECT  3.180 -0.210 3.640 0.210 ;
        RECT  2.920 -0.210 3.180 0.640 ;
        RECT  2.440 -0.210 2.920 0.210 ;
        RECT  2.220 -0.210 2.440 0.665 ;
        RECT  1.720 -0.210 2.220 0.210 ;
        RECT  1.500 -0.210 1.720 0.665 ;
        RECT  1.000 -0.210 1.500 0.210 ;
        RECT  0.780 -0.210 1.000 0.665 ;
        RECT  0.230 -0.210 0.780 0.210 ;
        RECT  0.090 -0.210 0.230 0.885 ;
        RECT  0.000 -0.210 0.090 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  21.670 2.310 21.840 2.730 ;
        RECT  21.540 1.655 21.670 2.730 ;
        RECT  20.965 2.310 21.540 2.730 ;
        RECT  20.795 1.665 20.965 2.730 ;
        RECT  20.245 2.310 20.795 2.730 ;
        RECT  20.075 1.665 20.245 2.730 ;
        RECT  19.525 2.310 20.075 2.730 ;
        RECT  19.355 1.665 19.525 2.730 ;
        RECT  18.805 2.310 19.355 2.730 ;
        RECT  18.635 1.665 18.805 2.730 ;
        RECT  18.130 2.310 18.635 2.730 ;
        RECT  17.870 1.830 18.130 2.730 ;
        RECT  17.410 2.310 17.870 2.730 ;
        RECT  17.150 2.035 17.410 2.730 ;
        RECT  16.190 2.310 17.150 2.730 ;
        RECT  15.930 1.875 16.190 2.730 ;
        RECT  15.260 2.310 15.930 2.730 ;
        RECT  15.000 2.130 15.260 2.730 ;
        RECT  14.520 2.310 15.000 2.730 ;
        RECT  14.260 2.130 14.520 2.730 ;
        RECT  13.760 2.310 14.260 2.730 ;
        RECT  13.500 2.130 13.760 2.730 ;
        RECT  13.005 2.310 13.500 2.730 ;
        RECT  12.745 2.130 13.005 2.730 ;
        RECT  12.240 2.310 12.745 2.730 ;
        RECT  11.980 2.130 12.240 2.730 ;
        RECT  11.360 2.310 11.980 2.730 ;
        RECT  11.100 2.220 11.360 2.730 ;
        RECT  8.640 2.310 11.100 2.730 ;
        RECT  8.380 2.220 8.640 2.730 ;
        RECT  7.880 2.310 8.380 2.730 ;
        RECT  7.620 2.220 7.880 2.730 ;
        RECT  7.020 2.310 7.620 2.730 ;
        RECT  6.760 2.220 7.020 2.730 ;
        RECT  5.870 2.310 6.760 2.730 ;
        RECT  5.610 2.055 5.870 2.730 ;
        RECT  4.610 2.310 5.610 2.730 ;
        RECT  4.350 2.055 4.610 2.730 ;
        RECT  3.855 2.310 4.350 2.730 ;
        RECT  3.685 1.665 3.855 2.730 ;
        RECT  3.135 2.310 3.685 2.730 ;
        RECT  2.965 1.665 3.135 2.730 ;
        RECT  2.415 2.310 2.965 2.730 ;
        RECT  2.240 1.655 2.415 2.730 ;
        RECT  1.695 2.310 2.240 2.730 ;
        RECT  1.520 1.655 1.695 2.730 ;
        RECT  0.975 2.310 1.520 2.730 ;
        RECT  0.800 1.655 0.975 2.730 ;
        RECT  0.230 2.310 0.800 2.730 ;
        RECT  0.100 1.655 0.230 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 21.840 2.520 ;
        LAYER M1 ;
        RECT  18.890 1.060 20.900 1.180 ;
        RECT  18.770 0.745 18.890 1.525 ;
        RECT  18.445 0.745 18.770 0.865 ;
        RECT  18.420 1.405 18.770 1.525 ;
        RECT  17.460 1.050 18.545 1.220 ;
        RECT  18.275 0.435 18.445 0.865 ;
        RECT  18.300 1.405 18.420 2.055 ;
        RECT  17.700 1.530 18.300 1.650 ;
        RECT  17.720 0.745 18.275 0.865 ;
        RECT  17.700 0.410 17.720 0.865 ;
        RECT  17.580 0.370 17.700 0.865 ;
        RECT  17.580 1.530 17.700 2.055 ;
        RECT  17.340 0.750 17.460 1.650 ;
        RECT  15.595 0.750 17.340 0.870 ;
        RECT  16.730 1.530 17.340 1.650 ;
        RECT  17.070 0.990 17.190 1.395 ;
        RECT  15.165 0.990 17.070 1.110 ;
        RECT  15.765 0.510 16.790 0.630 ;
        RECT  16.610 1.530 16.730 2.080 ;
        RECT  15.165 1.290 16.680 1.410 ;
        RECT  15.785 1.530 16.610 1.650 ;
        RECT  15.615 1.530 15.785 1.710 ;
        RECT  15.425 0.385 15.595 0.870 ;
        RECT  15.045 0.510 15.165 1.110 ;
        RECT  15.045 1.290 15.165 1.760 ;
        RECT  11.040 0.510 15.045 0.630 ;
        RECT  11.610 1.640 15.045 1.760 ;
        RECT  12.240 1.040 14.295 1.210 ;
        RECT  12.100 0.760 12.240 1.520 ;
        RECT  11.600 0.760 12.100 0.905 ;
        RECT  11.600 1.400 12.100 1.520 ;
        RECT  11.365 1.080 11.975 1.200 ;
        RECT  11.490 1.640 11.610 1.860 ;
        RECT  9.370 1.740 11.490 1.860 ;
        RECT  11.245 1.080 11.365 1.620 ;
        RECT  9.610 1.500 11.245 1.620 ;
        RECT  10.950 0.455 11.040 1.030 ;
        RECT  10.920 0.455 10.950 1.380 ;
        RECT  10.690 0.910 10.920 1.380 ;
        RECT  10.310 0.910 10.690 1.030 ;
        RECT  9.790 0.900 10.310 1.030 ;
        RECT  9.610 0.465 9.755 0.635 ;
        RECT  9.490 0.465 9.610 1.620 ;
        RECT  9.030 0.920 9.490 1.040 ;
        RECT  9.250 0.380 9.370 0.640 ;
        RECT  9.250 1.160 9.370 1.860 ;
        RECT  8.740 0.380 9.250 0.500 ;
        RECT  8.740 1.160 9.250 1.280 ;
        RECT  9.010 1.400 9.130 1.855 ;
        RECT  8.910 0.620 9.030 1.040 ;
        RECT  8.420 1.400 9.010 1.520 ;
        RECT  8.860 0.620 8.910 0.790 ;
        RECT  8.620 0.380 8.740 1.280 ;
        RECT  8.610 0.380 8.620 0.640 ;
        RECT  7.540 0.520 8.610 0.640 ;
        RECT  8.420 0.760 8.500 0.880 ;
        RECT  8.300 0.760 8.420 1.520 ;
        RECT  8.240 0.760 8.300 0.880 ;
        RECT  8.000 1.400 8.300 1.520 ;
        RECT  7.925 1.030 8.095 1.235 ;
        RECT  7.540 1.030 7.925 1.150 ;
        RECT  7.420 0.520 7.540 1.540 ;
        RECT  7.190 1.420 7.420 1.540 ;
        RECT  6.705 0.760 6.810 0.880 ;
        RECT  6.560 0.760 6.705 1.590 ;
        RECT  6.550 0.760 6.560 1.365 ;
        RECT  5.880 1.245 6.550 1.365 ;
        RECT  6.070 0.625 6.190 0.885 ;
        RECT  6.035 1.805 6.190 2.150 ;
        RECT  4.450 0.765 6.070 0.885 ;
        RECT  5.175 1.805 6.035 1.925 ;
        RECT  4.850 0.520 5.900 0.640 ;
        RECT  5.005 1.805 5.175 2.010 ;
        RECT  4.450 1.805 5.005 1.925 ;
        RECT  4.330 0.765 4.450 1.925 ;
        RECT  3.285 1.045 4.330 1.215 ;
        RECT  4.070 0.370 4.190 0.890 ;
        RECT  4.070 1.355 4.190 2.050 ;
        RECT  3.470 0.770 4.070 0.890 ;
        RECT  3.470 1.355 4.070 1.475 ;
        RECT  3.350 0.370 3.470 0.890 ;
        RECT  3.325 1.355 3.470 2.050 ;
        RECT  3.050 0.770 3.350 0.890 ;
        RECT  3.050 1.355 3.325 1.475 ;
        RECT  2.930 0.770 3.050 1.475 ;
        RECT  0.810 1.050 2.930 1.170 ;
    END
END BENCX4AD
MACRO BMXIX2AD
    CLASS CORE ;
    FOREIGN BMXIX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.625 1.910 5.885 2.170 ;
        END
        AntennaGateArea 0.1469 ;
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.210 0.980 4.410 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END S
    PIN PPN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.625 0.665 6.650 1.745 ;
        RECT  6.595 0.405 6.625 1.745 ;
        RECT  6.480 0.405 6.595 2.005 ;
        RECT  6.455 0.405 6.480 0.835 ;
        RECT  6.425 1.575 6.480 2.005 ;
        END
        AntennaDiffArea 0.373 ;
    END PPN
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.630 0.865 3.850 1.310 ;
        END
        AntennaGateArea 0.1468 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.400 0.860 1.520 2.090 ;
        RECT  1.260 1.970 1.400 2.090 ;
        RECT  1.000 1.970 1.260 2.190 ;
        RECT  0.490 1.970 1.000 2.090 ;
        RECT  0.430 1.160 0.490 2.090 ;
        RECT  0.350 1.020 0.430 2.090 ;
        RECT  0.310 1.020 0.350 1.280 ;
        END
        AntennaGateArea 0.1466 ;
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.615 1.040 0.770 1.455 ;
        END
        AntennaGateArea 0.1629 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.240 -0.210 6.720 0.210 ;
        RECT  5.980 -0.210 6.240 0.310 ;
        RECT  3.960 -0.210 5.980 0.210 ;
        RECT  3.700 -0.210 3.960 0.310 ;
        RECT  0.550 -0.210 3.700 0.210 ;
        RECT  0.290 -0.210 0.550 0.310 ;
        RECT  0.000 -0.210 0.290 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.250 2.310 6.720 2.730 ;
        RECT  6.050 1.565 6.250 2.730 ;
        RECT  3.945 2.310 6.050 2.730 ;
        RECT  3.685 2.210 3.945 2.730 ;
        RECT  0.550 2.310 3.685 2.730 ;
        RECT  0.290 2.210 0.550 2.730 ;
        RECT  0.000 2.310 0.290 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.720 2.520 ;
        LAYER M1 ;
        RECT  6.155 1.000 6.345 1.260 ;
        RECT  6.035 0.450 6.155 1.260 ;
        RECT  5.850 0.450 6.035 0.570 ;
        RECT  5.810 0.695 5.915 1.430 ;
        RECT  5.730 0.385 5.850 0.570 ;
        RECT  5.795 0.695 5.810 1.705 ;
        RECT  5.730 0.695 5.795 0.865 ;
        RECT  5.640 1.170 5.795 1.705 ;
        RECT  5.125 0.385 5.730 0.505 ;
        RECT  5.570 1.170 5.640 1.465 ;
        RECT  5.365 0.625 5.510 0.795 ;
        RECT  5.245 0.625 5.365 2.090 ;
        RECT  3.500 1.970 5.245 2.090 ;
        RECT  5.005 0.385 5.125 1.730 ;
        RECT  4.885 1.470 5.005 1.730 ;
        RECT  4.665 0.540 4.765 0.800 ;
        RECT  4.545 0.430 4.665 1.790 ;
        RECT  3.510 0.430 4.545 0.550 ;
        RECT  4.520 1.530 4.545 1.790 ;
        RECT  4.090 0.695 4.390 0.815 ;
        RECT  4.090 1.590 4.305 1.850 ;
        RECT  3.970 0.695 4.090 1.850 ;
        RECT  3.180 1.730 3.970 1.850 ;
        RECT  3.420 1.430 3.700 1.550 ;
        RECT  3.385 0.380 3.510 0.550 ;
        RECT  3.420 0.690 3.510 0.950 ;
        RECT  3.380 1.970 3.500 2.140 ;
        RECT  3.300 0.690 3.420 1.550 ;
        RECT  2.840 0.380 3.385 0.500 ;
        RECT  1.810 2.020 3.380 2.140 ;
        RECT  3.060 0.650 3.180 1.900 ;
        RECT  3.010 0.650 3.060 0.820 ;
        RECT  2.085 1.780 3.060 1.900 ;
        RECT  2.840 1.490 2.915 1.660 ;
        RECT  2.720 0.380 2.840 1.660 ;
        RECT  2.675 0.585 2.720 0.845 ;
        RECT  2.435 1.540 2.600 1.660 ;
        RECT  2.315 0.380 2.435 1.660 ;
        RECT  1.280 0.380 2.315 0.500 ;
        RECT  2.085 0.620 2.140 0.740 ;
        RECT  1.965 0.620 2.085 1.900 ;
        RECT  1.880 0.620 1.965 0.740 ;
        RECT  1.760 1.720 1.810 2.140 ;
        RECT  1.690 0.620 1.760 2.140 ;
        RECT  1.640 0.620 1.690 1.840 ;
        RECT  1.480 0.620 1.640 0.740 ;
        RECT  1.160 0.380 1.280 1.780 ;
        RECT  0.730 0.540 1.160 0.660 ;
        RECT  0.730 1.660 1.160 1.780 ;
        RECT  0.920 0.780 1.040 1.255 ;
        RECT  0.265 0.780 0.920 0.900 ;
        RECT  0.190 0.735 0.265 0.905 ;
        RECT  0.190 1.385 0.230 1.645 ;
        RECT  0.070 0.735 0.190 1.645 ;
    END
END BMXIX2AD
MACRO BMXIX4AD
    CLASS CORE ;
    FOREIGN BMXIX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.690 1.905 8.950 2.190 ;
        END
        AntennaGateArea 0.2734 ;
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.415 1.025 6.460 1.195 ;
        RECT  6.185 1.025 6.415 1.330 ;
        RECT  6.030 1.025 6.185 1.195 ;
        END
        AntennaGateArea 0.324 ;
    END S
    PIN PPN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.635 0.715 9.730 1.515 ;
        RECT  9.590 0.375 9.635 2.045 ;
        RECT  9.465 0.375 9.590 0.850 ;
        RECT  9.465 1.385 9.590 2.045 ;
        END
        AntennaDiffArea 0.422 ;
    END PPN
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 1.470 6.135 1.610 ;
        RECT  5.730 1.100 5.850 1.610 ;
        RECT  5.590 1.100 5.730 1.220 ;
        END
        AntennaGateArea 0.2734 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 0.880 1.990 1.955 ;
        RECT  1.635 1.835 1.870 1.955 ;
        RECT  1.515 1.835 1.635 2.190 ;
        RECT  0.490 1.835 1.515 1.955 ;
        RECT  0.350 1.005 0.490 1.955 ;
        END
        AntennaGateArea 0.2745 ;
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 1.015 1.170 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.970 -0.210 10.080 0.210 ;
        RECT  9.850 -0.210 9.970 0.595 ;
        RECT  9.250 -0.210 9.850 0.210 ;
        RECT  8.990 -0.210 9.250 0.310 ;
        RECT  6.855 -0.210 8.990 0.210 ;
        RECT  6.595 -0.210 6.855 0.310 ;
        RECT  5.950 -0.210 6.595 0.210 ;
        RECT  5.780 -0.210 5.950 0.310 ;
        RECT  1.460 -0.210 5.780 0.210 ;
        RECT  1.200 -0.210 1.460 0.400 ;
        RECT  0.710 -0.210 1.200 0.210 ;
        RECT  0.530 -0.210 0.710 0.515 ;
        RECT  0.000 -0.210 0.530 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.995 2.310 10.080 2.730 ;
        RECT  9.825 1.725 9.995 2.730 ;
        RECT  9.275 2.310 9.825 2.730 ;
        RECT  9.105 1.475 9.275 2.730 ;
        RECT  6.795 2.310 9.105 2.730 ;
        RECT  6.535 2.210 6.795 2.730 ;
        RECT  5.935 2.310 6.535 2.730 ;
        RECT  5.675 2.210 5.935 2.730 ;
        RECT  1.375 2.310 5.675 2.730 ;
        RECT  1.115 2.075 1.375 2.730 ;
        RECT  0.620 2.310 1.115 2.730 ;
        RECT  0.360 2.080 0.620 2.730 ;
        RECT  0.000 2.310 0.360 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.080 2.520 ;
        LAYER M1 ;
        RECT  9.340 0.985 9.460 1.245 ;
        RECT  9.205 0.985 9.340 1.105 ;
        RECT  9.085 0.495 9.205 1.105 ;
        RECT  8.420 0.495 9.085 0.615 ;
        RECT  8.885 0.735 8.920 0.905 ;
        RECT  8.750 0.735 8.885 1.785 ;
        RECT  8.710 1.210 8.750 1.785 ;
        RECT  8.540 1.210 8.710 1.470 ;
        RECT  8.300 0.380 8.420 1.900 ;
        RECT  7.795 0.380 8.300 0.500 ;
        RECT  8.250 1.470 8.300 1.900 ;
        RECT  8.035 0.675 8.180 1.035 ;
        RECT  8.010 0.675 8.035 2.090 ;
        RECT  7.915 0.915 8.010 2.090 ;
        RECT  5.570 1.970 7.915 2.090 ;
        RECT  7.675 0.380 7.795 0.775 ;
        RECT  7.555 0.380 7.675 1.850 ;
        RECT  6.985 1.730 7.555 1.850 ;
        RECT  7.315 0.430 7.435 1.610 ;
        RECT  5.650 0.430 7.315 0.550 ;
        RECT  7.125 1.490 7.315 1.610 ;
        RECT  6.985 0.670 7.145 0.790 ;
        RECT  6.835 0.670 6.985 1.850 ;
        RECT  6.585 0.745 6.705 1.850 ;
        RECT  6.165 0.745 6.585 0.865 ;
        RECT  5.320 1.730 6.585 1.850 ;
        RECT  5.540 0.695 5.710 0.980 ;
        RECT  5.530 0.380 5.650 0.550 ;
        RECT  5.440 1.410 5.600 1.530 ;
        RECT  5.450 1.970 5.570 2.140 ;
        RECT  5.440 0.860 5.540 0.980 ;
        RECT  4.960 0.380 5.530 0.500 ;
        RECT  2.255 2.020 5.450 2.140 ;
        RECT  5.320 0.860 5.440 1.530 ;
        RECT  5.200 0.620 5.415 0.740 ;
        RECT  5.200 1.730 5.320 1.900 ;
        RECT  5.080 0.620 5.200 1.900 ;
        RECT  3.770 1.780 5.080 1.900 ;
        RECT  4.840 0.380 4.960 1.660 ;
        RECT  4.170 1.540 4.840 1.660 ;
        RECT  4.480 0.380 4.600 1.420 ;
        RECT  3.425 0.380 4.480 0.500 ;
        RECT  4.320 1.300 4.480 1.420 ;
        RECT  4.170 0.620 4.310 0.740 ;
        RECT  4.050 0.620 4.170 1.660 ;
        RECT  3.940 1.540 4.050 1.660 ;
        RECT  3.770 0.620 3.930 0.740 ;
        RECT  3.650 0.620 3.770 1.900 ;
        RECT  2.640 1.780 3.650 1.900 ;
        RECT  3.290 0.380 3.425 1.660 ;
        RECT  1.925 0.380 3.290 0.500 ;
        RECT  3.165 1.540 3.290 1.660 ;
        RECT  2.255 0.620 3.120 0.740 ;
        RECT  2.610 0.860 2.740 0.980 ;
        RECT  2.610 1.715 2.640 1.900 ;
        RECT  2.470 0.860 2.610 1.900 ;
        RECT  2.135 0.620 2.255 2.140 ;
        RECT  2.095 0.620 2.135 0.740 ;
        RECT  1.805 0.380 1.925 0.730 ;
        RECT  1.750 0.520 1.805 0.730 ;
        RECT  1.630 0.520 1.750 1.715 ;
        RECT  1.055 0.520 1.630 0.640 ;
        RECT  1.580 1.515 1.630 1.715 ;
        RECT  0.755 1.515 1.580 1.635 ;
        RECT  1.390 0.760 1.510 1.210 ;
        RECT  0.270 0.760 1.390 0.880 ;
        RECT  0.885 0.435 1.055 0.640 ;
        RECT  0.230 0.605 0.270 0.880 ;
        RECT  0.110 0.605 0.230 1.670 ;
    END
END BMXIX4AD
MACRO BMXX2AD
    CLASS CORE ;
    FOREIGN BMXX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.695 1.875 6.795 2.135 ;
        RECT  6.415 1.875 6.695 2.170 ;
        RECT  6.185 2.030 6.415 2.170 ;
        END
        AntennaGateArea 0.1821 ;
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.990 0.915 4.225 1.375 ;
        END
        AntennaGateArea 0.1397 ;
    END S
    PIN PP
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.360 0.375 7.490 2.030 ;
        RECT  7.330 0.375 7.360 0.895 ;
        RECT  7.330 1.380 7.360 2.030 ;
        END
        AntennaDiffArea 0.373 ;
    END PP
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.690 0.785 3.850 1.305 ;
        RECT  3.665 0.910 3.690 1.305 ;
        END
        AntennaGateArea 0.1178 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.465 0.930 1.585 2.045 ;
        RECT  1.350 1.925 1.465 2.045 ;
        RECT  1.090 1.925 1.350 2.180 ;
        RECT  0.490 1.925 1.090 2.045 ;
        RECT  0.470 1.425 0.490 2.045 ;
        RECT  0.350 1.120 0.470 2.045 ;
        END
        AntennaGateArea 0.1173 ;
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.665 0.910 0.815 1.330 ;
        RECT  0.585 0.910 0.665 1.050 ;
        END
        AntennaGateArea 0.1403 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.090 -0.210 7.560 0.210 ;
        RECT  6.830 -0.210 7.090 0.265 ;
        RECT  5.245 -0.210 6.830 0.210 ;
        RECT  4.985 -0.210 5.245 0.255 ;
        RECT  4.075 -0.210 4.985 0.210 ;
        RECT  3.815 -0.210 4.075 0.260 ;
        RECT  0.660 -0.210 3.815 0.210 ;
        RECT  0.490 -0.210 0.660 0.550 ;
        RECT  0.000 -0.210 0.490 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.115 2.310 7.560 2.730 ;
        RECT  6.955 1.520 7.115 2.730 ;
        RECT  5.265 2.310 6.955 2.730 ;
        RECT  5.005 1.895 5.265 2.730 ;
        RECT  4.025 2.310 5.005 2.730 ;
        RECT  3.765 2.210 4.025 2.730 ;
        RECT  0.635 2.310 3.765 2.730 ;
        RECT  0.375 2.190 0.635 2.730 ;
        RECT  0.000 2.310 0.375 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  7.175 1.000 7.240 1.260 ;
        RECT  7.055 0.385 7.175 1.260 ;
        RECT  5.955 0.385 7.055 0.505 ;
        RECT  6.710 0.625 6.850 0.745 ;
        RECT  6.550 1.560 6.745 1.685 ;
        RECT  6.590 0.625 6.710 1.285 ;
        RECT  6.550 1.085 6.590 1.285 ;
        RECT  6.430 1.085 6.550 1.685 ;
        RECT  6.275 0.625 6.465 0.795 ;
        RECT  6.155 0.625 6.275 1.775 ;
        RECT  4.860 1.655 6.155 1.775 ;
        RECT  5.835 0.385 5.955 1.535 ;
        RECT  5.770 1.365 5.835 1.535 ;
        RECT  5.475 0.545 5.595 1.525 ;
        RECT  5.420 0.545 5.475 0.715 ;
        RECT  5.410 1.355 5.475 1.525 ;
        RECT  5.235 0.985 5.355 1.245 ;
        RECT  5.115 0.380 5.235 1.245 ;
        RECT  2.820 0.380 5.115 0.500 ;
        RECT  4.690 0.630 4.860 1.775 ;
        RECT  4.595 0.630 4.690 0.750 ;
        RECT  4.545 2.070 4.675 2.190 ;
        RECT  4.415 1.970 4.545 2.190 ;
        RECT  4.355 0.670 4.475 1.805 ;
        RECT  3.660 1.970 4.415 2.090 ;
        RECT  4.215 0.670 4.355 0.790 ;
        RECT  3.435 1.685 4.355 1.805 ;
        RECT  3.465 1.435 3.730 1.555 ;
        RECT  3.550 1.970 3.660 2.140 ;
        RECT  3.465 0.670 3.565 0.840 ;
        RECT  1.825 2.020 3.550 2.140 ;
        RECT  3.345 0.670 3.465 1.555 ;
        RECT  3.225 1.685 3.435 1.900 ;
        RECT  3.105 0.650 3.225 1.900 ;
        RECT  3.045 0.650 3.105 0.820 ;
        RECT  2.160 1.780 3.105 1.900 ;
        RECT  2.865 1.135 2.985 1.660 ;
        RECT  2.820 1.135 2.865 1.255 ;
        RECT  2.700 0.380 2.820 1.255 ;
        RECT  2.440 1.430 2.685 1.550 ;
        RECT  2.320 0.380 2.440 1.550 ;
        RECT  1.345 0.380 2.320 0.500 ;
        RECT  2.035 0.645 2.160 1.900 ;
        RECT  1.945 0.645 2.035 0.815 ;
        RECT  1.705 0.660 1.825 2.140 ;
        RECT  1.515 0.660 1.705 0.780 ;
        RECT  1.225 0.380 1.345 1.805 ;
        RECT  0.825 0.380 1.225 0.500 ;
        RECT  0.775 1.635 1.225 1.805 ;
        RECT  0.985 0.670 1.105 1.350 ;
        RECT  0.255 0.670 0.985 0.790 ;
        RECT  0.230 0.670 0.255 0.865 ;
        RECT  0.110 0.670 0.230 1.805 ;
        RECT  0.085 0.670 0.110 0.865 ;
    END
END BMXX2AD
MACRO BMXX4AD
    CLASS CORE ;
    FOREIGN BMXX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.295 2.030 8.685 2.180 ;
        END
        AntennaGateArea 0.3706 ;
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.225 0.950 4.455 1.330 ;
        END
        AntennaGateArea 0.2788 ;
    END S
    PIN PP
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.355 0.660 9.450 1.515 ;
        RECT  9.310 0.420 9.355 1.995 ;
        RECT  9.185 0.420 9.310 0.850 ;
        RECT  9.185 1.380 9.310 1.995 ;
        END
        AntennaDiffArea 0.419 ;
    END PP
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.470 4.175 1.610 ;
        RECT  3.940 1.105 4.060 1.610 ;
        RECT  3.845 1.105 3.940 1.300 ;
        END
        AntennaGateArea 0.1874 ;
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.160 1.265 ;
        RECT  0.910 1.005 1.050 1.375 ;
        END
        AntennaGateArea 0.1873 ;
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.015 0.785 1.375 ;
        RECT  0.360 1.015 0.630 1.275 ;
        END
        AntennaGateArea 0.278 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.690 -0.210 9.800 0.210 ;
        RECT  9.570 -0.210 9.690 0.805 ;
        RECT  9.020 -0.210 9.570 0.210 ;
        RECT  8.760 -0.210 9.020 0.260 ;
        RECT  6.590 -0.210 8.760 0.210 ;
        RECT  6.330 -0.210 6.590 0.260 ;
        RECT  5.830 -0.210 6.330 0.210 ;
        RECT  5.570 -0.210 5.830 0.310 ;
        RECT  5.040 -0.210 5.570 0.210 ;
        RECT  4.780 -0.210 5.040 0.310 ;
        RECT  4.245 -0.210 4.780 0.210 ;
        RECT  3.985 -0.210 4.245 0.310 ;
        RECT  1.050 -0.210 3.985 0.210 ;
        RECT  0.790 -0.210 1.050 0.325 ;
        RECT  0.265 -0.210 0.790 0.210 ;
        RECT  0.095 -0.210 0.265 0.585 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.690 2.310 9.800 2.730 ;
        RECT  9.570 1.675 9.690 2.730 ;
        RECT  8.970 2.310 9.570 2.730 ;
        RECT  8.850 1.435 8.970 2.730 ;
        RECT  6.460 2.310 8.850 2.730 ;
        RECT  6.200 2.190 6.460 2.730 ;
        RECT  5.690 2.310 6.200 2.730 ;
        RECT  5.430 2.190 5.690 2.730 ;
        RECT  4.930 2.310 5.430 2.730 ;
        RECT  4.670 2.220 4.930 2.730 ;
        RECT  4.170 2.310 4.670 2.730 ;
        RECT  3.910 2.220 4.170 2.730 ;
        RECT  1.025 2.310 3.910 2.730 ;
        RECT  0.855 1.555 1.025 2.730 ;
        RECT  0.305 2.310 0.855 2.730 ;
        RECT  0.135 1.735 0.305 2.730 ;
        RECT  0.000 2.310 0.135 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.800 2.520 ;
        LAYER M1 ;
        RECT  9.060 0.985 9.180 1.245 ;
        RECT  8.970 0.985 9.060 1.120 ;
        RECT  8.850 0.380 8.970 1.120 ;
        RECT  8.180 0.380 8.850 0.500 ;
        RECT  8.530 0.630 8.640 0.750 ;
        RECT  8.530 1.465 8.595 1.895 ;
        RECT  8.380 0.630 8.530 1.895 ;
        RECT  8.235 1.120 8.380 1.380 ;
        RECT  8.110 0.380 8.180 1.000 ;
        RECT  8.060 0.380 8.110 1.890 ;
        RECT  7.510 0.380 8.060 0.500 ;
        RECT  7.990 0.865 8.060 1.890 ;
        RECT  7.800 0.620 7.940 0.740 ;
        RECT  7.750 0.620 7.800 1.200 ;
        RECT  7.680 0.620 7.750 2.055 ;
        RECT  7.630 1.080 7.680 2.055 ;
        RECT  5.405 1.935 7.630 2.055 ;
        RECT  7.390 0.380 7.510 1.815 ;
        RECT  6.670 1.695 7.390 1.815 ;
        RECT  7.030 0.380 7.165 1.575 ;
        RECT  6.430 0.380 7.030 0.500 ;
        RECT  6.840 1.455 7.030 1.575 ;
        RECT  6.670 0.620 6.860 0.740 ;
        RECT  6.550 0.620 6.670 1.815 ;
        RECT  6.310 0.380 6.430 1.745 ;
        RECT  6.165 0.685 6.310 0.805 ;
        RECT  6.025 1.625 6.310 1.745 ;
        RECT  5.995 0.565 6.165 0.805 ;
        RECT  5.790 1.070 6.145 1.240 ;
        RECT  5.855 1.625 6.025 1.795 ;
        RECT  5.670 0.430 5.790 1.240 ;
        RECT  3.840 0.430 5.670 0.550 ;
        RECT  5.275 0.670 5.405 2.055 ;
        RECT  5.235 0.670 5.275 0.840 ;
        RECT  5.120 1.535 5.275 2.055 ;
        RECT  5.000 1.060 5.145 1.230 ;
        RECT  4.880 1.060 5.000 2.100 ;
        RECT  3.700 1.980 4.880 2.100 ;
        RECT  4.575 0.705 4.695 1.860 ;
        RECT  4.365 0.705 4.575 0.825 ;
        RECT  3.450 1.740 4.575 1.860 ;
        RECT  3.725 0.705 3.895 0.985 ;
        RECT  3.720 0.380 3.840 0.550 ;
        RECT  3.630 1.500 3.820 1.620 ;
        RECT  3.630 0.865 3.725 0.985 ;
        RECT  3.150 0.380 3.720 0.500 ;
        RECT  3.580 1.980 3.700 2.140 ;
        RECT  3.510 0.865 3.630 1.620 ;
        RECT  3.390 0.620 3.580 0.740 ;
        RECT  1.640 2.020 3.580 2.140 ;
        RECT  3.390 1.740 3.450 1.900 ;
        RECT  3.270 0.620 3.390 1.900 ;
        RECT  2.325 1.780 3.270 1.900 ;
        RECT  3.085 0.380 3.150 1.335 ;
        RECT  3.030 0.380 3.085 1.660 ;
        RECT  2.965 1.215 3.030 1.660 ;
        RECT  2.825 1.540 2.965 1.660 ;
        RECT  2.705 0.380 2.790 1.065 ;
        RECT  2.670 0.380 2.705 1.660 ;
        RECT  1.735 0.380 2.670 0.500 ;
        RECT  2.585 0.945 2.670 1.660 ;
        RECT  2.445 1.540 2.585 1.660 ;
        RECT  2.380 0.645 2.465 0.815 ;
        RECT  2.325 0.645 2.380 1.345 ;
        RECT  2.260 0.645 2.325 1.900 ;
        RECT  2.205 1.225 2.260 1.900 ;
        RECT  1.880 1.780 2.205 1.900 ;
        RECT  1.985 0.640 2.140 0.760 ;
        RECT  1.865 0.640 1.985 1.380 ;
        RECT  1.760 1.640 1.880 1.900 ;
        RECT  1.640 1.260 1.865 1.380 ;
        RECT  1.565 0.355 1.735 0.785 ;
        RECT  1.400 1.015 1.690 1.135 ;
        RECT  1.520 1.260 1.640 2.140 ;
        RECT  1.005 0.445 1.565 0.565 ;
        RECT  1.280 0.705 1.400 1.635 ;
        RECT  1.215 0.705 1.280 0.875 ;
        RECT  1.240 1.375 1.280 1.635 ;
        RECT  0.885 0.445 1.005 0.825 ;
        RECT  0.625 0.705 0.885 0.825 ;
        RECT  0.495 1.495 0.665 1.940 ;
        RECT  0.455 0.375 0.625 0.825 ;
        RECT  0.210 1.495 0.495 1.615 ;
        RECT  0.210 0.705 0.455 0.825 ;
        RECT  0.090 0.705 0.210 1.615 ;
    END
END BMXX4AD
MACRO BUFX10AD
    CLASS CORE ;
    FOREIGN BUFX10AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.670 0.380 2.840 2.125 ;
        RECT  2.190 0.695 2.670 1.675 ;
        RECT  2.145 0.695 2.190 2.125 ;
        RECT  2.010 0.380 2.145 2.125 ;
        RECT  1.925 0.380 2.010 0.925 ;
        RECT  1.885 1.385 2.010 2.125 ;
        RECT  1.425 0.695 1.925 0.925 ;
        RECT  1.465 1.385 1.885 1.615 ;
        RECT  1.210 1.385 1.465 2.125 ;
        RECT  1.195 0.375 1.425 0.925 ;
        END
        AntennaDiffArea 1.217 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 1.020 0.505 1.280 ;
        RECT  0.215 1.020 0.310 1.375 ;
        RECT  0.070 1.135 0.215 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.525 -0.210 3.080 0.210 ;
        RECT  2.265 -0.210 2.525 0.500 ;
        RECT  1.805 -0.210 2.265 0.210 ;
        RECT  1.545 -0.210 1.805 0.500 ;
        RECT  1.040 -0.210 1.545 0.210 ;
        RECT  0.870 -0.210 1.040 0.815 ;
        RECT  0.320 -0.210 0.870 0.210 ;
        RECT  0.150 -0.210 0.320 0.835 ;
        RECT  0.000 -0.210 0.150 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 2.310 3.080 2.730 ;
        RECT  2.310 1.860 2.480 2.730 ;
        RECT  1.760 2.310 2.310 2.730 ;
        RECT  1.590 1.780 1.760 2.730 ;
        RECT  1.015 2.310 1.590 2.730 ;
        RECT  0.895 1.525 1.015 2.730 ;
        RECT  0.335 2.310 0.895 2.730 ;
        RECT  0.145 1.530 0.335 2.730 ;
        RECT  0.000 2.310 0.145 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  0.745 1.095 1.765 1.215 ;
        RECT  0.680 0.380 0.745 1.660 ;
        RECT  0.625 0.380 0.680 2.185 ;
        RECT  0.510 0.380 0.625 0.810 ;
        RECT  0.510 1.495 0.625 2.185 ;
    END
END BUFX10AD
MACRO BUFX12AD
    CLASS CORE ;
    FOREIGN BUFX12AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.995 0.375 3.165 2.110 ;
        RECT  2.965 0.540 2.995 2.110 ;
        RECT  2.480 0.540 2.965 1.725 ;
        RECT  2.450 0.540 2.480 2.115 ;
        RECT  2.290 0.360 2.450 2.115 ;
        RECT  2.250 0.360 2.290 0.900 ;
        RECT  2.240 1.360 2.290 2.115 ;
        RECT  1.750 0.540 2.250 0.900 ;
        RECT  1.725 1.360 2.240 1.725 ;
        RECT  1.530 0.360 1.750 0.900 ;
        RECT  1.555 1.360 1.725 2.115 ;
        END
        AntennaDiffArea 1.266 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.345 1.085 0.775 1.375 ;
        END
        AntennaGateArea 0.3878 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 -0.210 3.640 0.210 ;
        RECT  3.355 -0.210 3.525 0.800 ;
        RECT  2.850 -0.210 3.355 0.210 ;
        RECT  2.590 -0.210 2.850 0.420 ;
        RECT  2.130 -0.210 2.590 0.210 ;
        RECT  1.870 -0.210 2.130 0.420 ;
        RECT  1.365 -0.210 1.870 0.210 ;
        RECT  1.195 -0.210 1.365 0.840 ;
        RECT  0.645 -0.210 1.195 0.210 ;
        RECT  0.475 -0.210 0.645 0.680 ;
        RECT  0.000 -0.210 0.475 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.525 2.310 3.640 2.730 ;
        RECT  3.355 1.455 3.525 2.730 ;
        RECT  2.805 2.310 3.355 2.730 ;
        RECT  2.635 1.845 2.805 2.730 ;
        RECT  2.085 2.310 2.635 2.730 ;
        RECT  1.915 1.845 2.085 2.730 ;
        RECT  1.365 2.310 1.915 2.730 ;
        RECT  1.195 1.530 1.365 2.730 ;
        RECT  0.645 2.310 1.195 2.730 ;
        RECT  0.475 1.540 0.645 2.730 ;
        RECT  0.000 2.310 0.475 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  1.015 1.070 2.170 1.190 ;
        RECT  0.895 0.425 1.015 1.970 ;
        RECT  0.835 0.425 0.895 0.930 ;
        RECT  0.835 1.540 0.895 1.970 ;
        RECT  0.275 0.810 0.835 0.930 ;
        RECT  0.225 0.445 0.275 0.930 ;
        RECT  0.225 1.540 0.275 1.970 ;
        RECT  0.105 0.445 0.225 1.970 ;
    END
END BUFX12AD
MACRO BUFX14AD
    CLASS CORE ;
    FOREIGN BUFX14AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.785 0.420 3.955 0.920 ;
        RECT  3.785 1.310 3.955 2.120 ;
        RECT  3.310 0.560 3.785 0.920 ;
        RECT  3.310 1.310 3.785 1.765 ;
        RECT  3.250 0.560 3.310 1.765 ;
        RECT  3.050 0.375 3.250 2.130 ;
        RECT  2.570 0.560 3.050 1.765 ;
        RECT  2.540 0.560 2.570 0.920 ;
        RECT  2.550 1.380 2.570 1.765 ;
        RECT  2.300 1.380 2.550 2.130 ;
        RECT  2.320 0.405 2.540 0.920 ;
        RECT  1.820 0.560 2.320 0.920 ;
        RECT  1.795 1.380 2.300 1.765 ;
        RECT  1.570 0.400 1.820 0.920 ;
        RECT  1.625 1.380 1.795 2.115 ;
        END
        AntennaDiffArea 1.639 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.110 0.900 1.230 ;
        RECT  0.350 1.110 0.770 1.375 ;
        END
        AntennaGateArea 0.4539 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.640 -0.210 4.200 0.210 ;
        RECT  3.380 -0.210 3.640 0.440 ;
        RECT  2.920 -0.210 3.380 0.210 ;
        RECT  2.660 -0.210 2.920 0.440 ;
        RECT  2.200 -0.210 2.660 0.210 ;
        RECT  1.940 -0.210 2.200 0.440 ;
        RECT  1.435 -0.210 1.940 0.210 ;
        RECT  1.265 -0.210 1.435 0.820 ;
        RECT  0.715 -0.210 1.265 0.210 ;
        RECT  0.545 -0.210 0.715 0.735 ;
        RECT  0.000 -0.210 0.545 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.595 2.310 4.200 2.730 ;
        RECT  3.425 1.890 3.595 2.730 ;
        RECT  2.875 2.310 3.425 2.730 ;
        RECT  2.705 1.890 2.875 2.730 ;
        RECT  2.155 2.310 2.705 2.730 ;
        RECT  1.985 1.885 2.155 2.730 ;
        RECT  1.435 2.310 1.985 2.730 ;
        RECT  1.265 1.465 1.435 2.730 ;
        RECT  0.715 2.310 1.265 2.730 ;
        RECT  0.545 1.785 0.715 2.730 ;
        RECT  0.000 2.310 0.545 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  1.140 1.090 2.240 1.210 ;
        RECT  1.075 0.855 1.140 1.665 ;
        RECT  1.020 0.430 1.075 2.185 ;
        RECT  0.905 0.430 1.020 0.975 ;
        RECT  0.905 1.495 1.020 2.185 ;
        RECT  0.355 0.855 0.905 0.975 ;
        RECT  0.355 1.545 0.905 1.665 ;
        RECT  0.185 0.435 0.355 0.975 ;
        RECT  0.185 1.545 0.355 2.060 ;
    END
END BUFX14AD
MACRO BUFX16AD
    CLASS CORE ;
    FOREIGN BUFX16AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.685 0.380 3.855 0.920 ;
        RECT  3.685 1.380 3.855 2.075 ;
        RECT  3.590 0.510 3.685 0.920 ;
        RECT  3.590 1.380 3.685 1.880 ;
        RECT  3.135 0.510 3.590 1.880 ;
        RECT  2.965 0.390 3.135 2.085 ;
        RECT  2.850 0.510 2.965 1.880 ;
        RECT  2.440 0.510 2.850 0.920 ;
        RECT  2.415 1.380 2.850 1.880 ;
        RECT  2.220 0.405 2.440 0.920 ;
        RECT  2.245 1.380 2.415 2.115 ;
        RECT  1.695 1.380 2.245 1.880 ;
        RECT  1.720 0.510 2.220 0.920 ;
        RECT  1.470 0.400 1.720 0.920 ;
        RECT  1.525 1.380 1.695 2.115 ;
        END
        AntennaDiffArea 1.736 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.140 0.800 1.260 ;
        RECT  0.070 1.140 0.490 1.375 ;
        END
        AntennaGateArea 0.4869 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.245 -0.210 4.480 0.210 ;
        RECT  4.075 -0.210 4.245 0.825 ;
        RECT  3.540 -0.210 4.075 0.210 ;
        RECT  3.280 -0.210 3.540 0.390 ;
        RECT  2.820 -0.210 3.280 0.210 ;
        RECT  2.560 -0.210 2.820 0.390 ;
        RECT  2.100 -0.210 2.560 0.210 ;
        RECT  1.840 -0.210 2.100 0.390 ;
        RECT  1.335 -0.210 1.840 0.210 ;
        RECT  1.165 -0.210 1.335 0.830 ;
        RECT  0.615 -0.210 1.165 0.210 ;
        RECT  0.445 -0.210 0.615 0.745 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.245 2.310 4.480 2.730 ;
        RECT  4.075 1.480 4.245 2.730 ;
        RECT  3.495 2.310 4.075 2.730 ;
        RECT  3.325 2.010 3.495 2.730 ;
        RECT  2.775 2.310 3.325 2.730 ;
        RECT  2.605 2.015 2.775 2.730 ;
        RECT  2.055 2.310 2.605 2.730 ;
        RECT  1.885 2.010 2.055 2.730 ;
        RECT  1.335 2.310 1.885 2.730 ;
        RECT  1.165 1.490 1.335 2.730 ;
        RECT  0.615 2.310 1.165 2.730 ;
        RECT  0.445 1.755 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
        LAYER M1 ;
        RECT  1.040 1.090 2.660 1.210 ;
        RECT  0.975 0.420 1.040 1.615 ;
        RECT  0.920 0.420 0.975 2.185 ;
        RECT  0.805 0.420 0.920 1.000 ;
        RECT  0.805 1.495 0.920 2.185 ;
        RECT  0.255 0.880 0.805 1.000 ;
        RECT  0.255 1.495 0.805 1.615 ;
        RECT  0.085 0.425 0.255 1.000 ;
        RECT  0.085 1.495 0.255 2.185 ;
    END
END BUFX16AD
MACRO BUFX18AD
    CLASS CORE ;
    FOREIGN BUFX18AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.765 0.405 4.935 0.920 ;
        RECT  4.765 1.380 4.935 2.070 ;
        RECT  4.215 0.530 4.765 0.920 ;
        RECT  4.215 1.380 4.765 1.880 ;
        RECT  4.185 0.410 4.215 0.920 ;
        RECT  4.185 1.380 4.215 2.070 ;
        RECT  4.045 0.410 4.185 2.070 ;
        RECT  3.495 0.530 4.045 1.880 ;
        RECT  3.325 0.410 3.495 2.070 ;
        RECT  2.775 0.530 3.325 0.920 ;
        RECT  2.775 1.380 3.325 1.880 ;
        RECT  2.605 0.435 2.775 0.920 ;
        RECT  2.605 1.380 2.775 2.070 ;
        RECT  2.080 0.530 2.605 0.920 ;
        RECT  2.055 1.380 2.605 1.880 ;
        RECT  1.830 0.400 2.080 0.920 ;
        RECT  1.885 1.380 2.055 2.070 ;
        END
        AntennaDiffArea 2.061 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.120 1.060 1.240 ;
        RECT  0.070 1.120 0.490 1.375 ;
        END
        AntennaGateArea 0.584 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.620 -0.210 5.040 0.210 ;
        RECT  4.360 -0.210 4.620 0.400 ;
        RECT  3.900 -0.210 4.360 0.210 ;
        RECT  3.640 -0.210 3.900 0.400 ;
        RECT  3.180 -0.210 3.640 0.210 ;
        RECT  2.920 -0.210 3.180 0.400 ;
        RECT  2.460 -0.210 2.920 0.210 ;
        RECT  2.200 -0.210 2.460 0.400 ;
        RECT  1.695 -0.210 2.200 0.210 ;
        RECT  1.525 -0.210 1.695 0.890 ;
        RECT  0.975 -0.210 1.525 0.210 ;
        RECT  0.805 -0.210 0.975 0.755 ;
        RECT  0.255 -0.210 0.805 0.210 ;
        RECT  0.085 -0.210 0.255 0.860 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.575 2.310 5.040 2.730 ;
        RECT  4.405 2.005 4.575 2.730 ;
        RECT  3.855 2.310 4.405 2.730 ;
        RECT  3.685 2.005 3.855 2.730 ;
        RECT  3.135 2.310 3.685 2.730 ;
        RECT  2.965 2.005 3.135 2.730 ;
        RECT  2.415 2.310 2.965 2.730 ;
        RECT  2.245 2.000 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 1.465 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.735 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.505 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.040 2.520 ;
        LAYER M1 ;
        RECT  1.370 1.090 3.020 1.210 ;
        RECT  1.335 0.450 1.370 1.615 ;
        RECT  1.250 0.450 1.335 2.185 ;
        RECT  1.165 0.450 1.250 1.000 ;
        RECT  1.165 1.495 1.250 2.185 ;
        RECT  0.615 0.880 1.165 1.000 ;
        RECT  0.615 1.495 1.165 1.615 ;
        RECT  0.445 0.390 0.615 1.000 ;
        RECT  0.445 1.495 0.615 2.185 ;
    END
END BUFX18AD
MACRO BUFX20AD
    CLASS CORE ;
    FOREIGN BUFX20AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.765 0.405 4.935 0.920 ;
        RECT  4.765 1.380 4.935 2.070 ;
        RECT  4.215 0.520 4.765 0.920 ;
        RECT  4.215 1.380 4.765 1.980 ;
        RECT  4.185 0.410 4.215 0.920 ;
        RECT  4.185 1.380 4.215 2.070 ;
        RECT  4.045 0.410 4.185 2.070 ;
        RECT  3.495 0.520 4.045 1.980 ;
        RECT  3.325 0.410 3.495 2.070 ;
        RECT  2.775 0.520 3.325 0.920 ;
        RECT  2.775 1.380 3.325 1.980 ;
        RECT  2.605 0.435 2.775 0.920 ;
        RECT  2.605 1.380 2.775 2.070 ;
        RECT  2.080 0.520 2.605 0.920 ;
        RECT  2.055 1.380 2.605 1.980 ;
        RECT  1.830 0.400 2.080 0.920 ;
        RECT  1.885 1.380 2.055 2.070 ;
        END
        AntennaDiffArea 2.11 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.120 1.060 1.240 ;
        RECT  0.070 1.120 0.490 1.375 ;
        END
        AntennaGateArea 0.648 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.295 -0.210 5.600 0.210 ;
        RECT  5.125 -0.210 5.295 0.835 ;
        RECT  4.620 -0.210 5.125 0.210 ;
        RECT  4.360 -0.210 4.620 0.400 ;
        RECT  3.900 -0.210 4.360 0.210 ;
        RECT  3.640 -0.210 3.900 0.400 ;
        RECT  3.180 -0.210 3.640 0.210 ;
        RECT  2.920 -0.210 3.180 0.400 ;
        RECT  2.460 -0.210 2.920 0.210 ;
        RECT  2.200 -0.210 2.460 0.400 ;
        RECT  1.695 -0.210 2.200 0.210 ;
        RECT  1.525 -0.210 1.695 0.890 ;
        RECT  0.975 -0.210 1.525 0.210 ;
        RECT  0.805 -0.210 0.975 0.755 ;
        RECT  0.255 -0.210 0.805 0.210 ;
        RECT  0.085 -0.210 0.255 0.860 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.295 2.310 5.600 2.730 ;
        RECT  5.125 1.450 5.295 2.730 ;
        RECT  4.620 2.310 5.125 2.730 ;
        RECT  4.360 2.105 4.620 2.730 ;
        RECT  3.900 2.310 4.360 2.730 ;
        RECT  3.640 2.105 3.900 2.730 ;
        RECT  3.180 2.310 3.640 2.730 ;
        RECT  2.920 2.105 3.180 2.730 ;
        RECT  2.460 2.310 2.920 2.730 ;
        RECT  2.200 2.105 2.460 2.730 ;
        RECT  1.695 2.310 2.200 2.730 ;
        RECT  1.525 1.465 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.735 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.545 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  1.370 1.090 3.020 1.210 ;
        RECT  1.335 0.450 1.370 1.615 ;
        RECT  1.250 0.450 1.335 2.185 ;
        RECT  1.165 0.450 1.250 1.000 ;
        RECT  1.165 1.495 1.250 2.185 ;
        RECT  0.615 0.880 1.165 1.000 ;
        RECT  0.615 1.495 1.165 1.615 ;
        RECT  0.445 0.390 0.615 1.000 ;
        RECT  0.445 1.495 0.615 2.185 ;
    END
END BUFX20AD
MACRO BUFX2AD
    CLASS CORE ;
    FOREIGN BUFX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.365 1.050 2.035 ;
        RECT  0.880 0.365 0.910 0.885 ;
        RECT  0.880 1.515 0.910 2.035 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.065 0.375 1.235 ;
        RECT  0.070 1.065 0.210 1.375 ;
        END
        AntennaGateArea 0.0651 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.720 -0.210 1.120 0.210 ;
        RECT  0.460 -0.210 0.720 0.540 ;
        RECT  0.000 -0.210 0.460 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.675 2.310 1.120 2.730 ;
        RECT  0.505 1.780 0.675 2.730 ;
        RECT  0.000 2.310 0.505 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
        LAYER M1 ;
        RECT  0.625 0.690 0.745 1.615 ;
        RECT  0.085 0.690 0.625 0.860 ;
        RECT  0.255 1.495 0.625 1.615 ;
        RECT  0.085 1.495 0.255 1.665 ;
    END
END BUFX2AD
MACRO BUFX3AD
    CLASS CORE ;
    FOREIGN BUFX3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.605 1.050 1.940 ;
        RECT  0.810 0.605 0.910 0.865 ;
        RECT  0.810 1.420 0.910 1.940 ;
        END
        AntennaDiffArea 0.318 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.285 1.090 0.450 1.210 ;
        RECT  0.210 1.065 0.285 1.235 ;
        RECT  0.070 1.065 0.210 1.375 ;
        END
        AntennaGateArea 0.0984 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.300 -0.210 1.400 0.210 ;
        RECT  1.170 -0.210 1.300 0.810 ;
        RECT  0.620 -0.210 1.170 0.210 ;
        RECT  0.360 -0.210 0.620 0.240 ;
        RECT  0.000 -0.210 0.360 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.295 2.310 1.400 2.730 ;
        RECT  1.170 1.465 1.295 2.730 ;
        RECT  0.575 2.310 1.170 2.730 ;
        RECT  0.405 2.175 0.575 2.730 ;
        RECT  0.000 2.310 0.405 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.690 1.030 0.790 1.290 ;
        RECT  0.570 0.660 0.690 1.685 ;
        RECT  0.085 0.660 0.570 0.830 ;
        RECT  0.085 1.515 0.570 1.685 ;
    END
END BUFX3AD
MACRO BUFX4AD
    CLASS CORE ;
    FOREIGN BUFX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.345 0.825 1.475 1.560 ;
        RECT  1.065 0.825 1.345 0.955 ;
        RECT  1.075 1.400 1.345 1.560 ;
        RECT  0.895 1.400 1.075 2.055 ;
        RECT  0.895 0.400 1.065 0.955 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.490 1.375 ;
        END
        AntennaGateArea 0.1297 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.425 -0.210 1.680 0.210 ;
        RECT  1.255 -0.210 1.425 0.695 ;
        RECT  0.705 -0.210 1.255 0.210 ;
        RECT  0.535 -0.210 0.705 0.725 ;
        RECT  0.000 -0.210 0.535 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.425 2.310 1.680 2.730 ;
        RECT  1.255 1.735 1.425 2.730 ;
        RECT  0.705 2.310 1.255 2.730 ;
        RECT  0.535 1.735 0.705 2.730 ;
        RECT  0.000 2.310 0.535 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  0.775 1.105 1.220 1.225 ;
        RECT  0.655 1.105 0.775 1.615 ;
        RECT  0.305 1.495 0.655 1.615 ;
        RECT  0.230 1.495 0.305 1.925 ;
        RECT  0.230 0.510 0.295 0.730 ;
        RECT  0.110 0.510 0.230 1.925 ;
    END
END BUFX4AD
MACRO BUFX5AD
    CLASS CORE ;
    FOREIGN BUFX5AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.415 1.815 2.110 ;
        RECT  1.075 0.780 1.630 0.955 ;
        RECT  1.075 1.345 1.630 1.515 ;
        RECT  0.865 0.400 1.075 0.955 ;
        RECT  0.885 1.345 1.075 2.125 ;
        END
        AntennaDiffArea 0.656 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.975 0.525 1.375 ;
        END
        AntennaGateArea 0.161 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.395 -0.210 1.960 0.210 ;
        RECT  1.225 -0.210 1.395 0.635 ;
        RECT  0.680 -0.210 1.225 0.210 ;
        RECT  0.460 -0.210 0.680 0.795 ;
        RECT  0.000 -0.210 0.460 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.395 2.310 1.960 2.730 ;
        RECT  1.225 1.655 1.395 2.730 ;
        RECT  0.645 2.310 1.225 2.730 ;
        RECT  0.475 1.815 0.645 2.730 ;
        RECT  0.000 2.310 0.475 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  0.765 1.095 1.510 1.215 ;
        RECT  0.645 1.095 0.765 1.615 ;
        RECT  0.285 1.495 0.645 1.615 ;
        RECT  0.230 0.345 0.285 0.775 ;
        RECT  0.230 1.495 0.285 2.185 ;
        RECT  0.105 0.345 0.230 2.185 ;
    END
END BUFX5AD
MACRO BUFX6AD
    CLASS CORE ;
    FOREIGN BUFX6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.905 0.370 2.135 2.135 ;
        RECT  1.890 0.370 1.905 1.660 ;
        RECT  1.750 0.660 1.890 1.660 ;
        RECT  1.430 0.660 1.750 0.920 ;
        RECT  1.460 1.365 1.750 1.660 ;
        RECT  1.220 1.365 1.460 2.135 ;
        RECT  1.225 0.415 1.430 0.920 ;
        END
        AntennaDiffArea 0.795 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.105 0.795 1.225 ;
        RECT  0.070 1.105 0.210 1.375 ;
        END
        AntennaGateArea 0.1972 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.210 2.240 0.210 ;
        RECT  1.585 -0.210 1.765 0.535 ;
        RECT  1.035 -0.210 1.585 0.210 ;
        RECT  0.865 -0.210 1.035 0.725 ;
        RECT  0.270 -0.210 0.865 0.210 ;
        RECT  0.100 -0.210 0.270 0.875 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.775 2.310 2.240 2.730 ;
        RECT  1.605 1.845 1.775 2.730 ;
        RECT  1.040 2.310 1.605 2.730 ;
        RECT  0.840 1.585 1.040 2.730 ;
        RECT  0.270 2.310 0.840 2.730 ;
        RECT  0.100 1.545 0.270 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.095 1.080 1.580 1.200 ;
        RECT  0.930 0.850 1.095 1.465 ;
        RECT  0.630 0.850 0.930 0.970 ;
        RECT  0.650 1.345 0.930 1.465 ;
        RECT  0.460 1.345 0.650 1.895 ;
        RECT  0.460 0.660 0.630 0.970 ;
    END
END BUFX6AD
MACRO BUFX8AD
    CLASS CORE ;
    FOREIGN BUFX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.905 0.465 2.075 2.110 ;
        RECT  1.855 0.645 1.905 2.110 ;
        RECT  1.610 0.645 1.855 1.565 ;
        RECT  1.380 0.645 1.610 0.925 ;
        RECT  1.400 1.335 1.610 1.565 ;
        RECT  1.150 1.335 1.400 2.115 ;
        RECT  1.165 0.395 1.380 0.925 ;
        END
        AntennaDiffArea 0.854 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.040 0.710 1.375 ;
        END
        AntennaGateArea 0.258 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 -0.210 2.520 0.210 ;
        RECT  2.265 -0.210 2.435 0.825 ;
        RECT  1.715 -0.210 2.265 0.210 ;
        RECT  1.545 -0.210 1.715 0.525 ;
        RECT  0.995 -0.210 1.545 0.210 ;
        RECT  0.825 -0.210 0.995 0.610 ;
        RECT  0.265 -0.210 0.825 0.210 ;
        RECT  0.095 -0.210 0.265 0.835 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 2.310 2.520 2.730 ;
        RECT  2.265 1.450 2.435 2.730 ;
        RECT  1.705 2.310 2.265 2.730 ;
        RECT  1.535 1.735 1.705 2.730 ;
        RECT  0.985 2.310 1.535 2.730 ;
        RECT  0.815 1.790 0.985 2.730 ;
        RECT  0.265 2.310 0.815 2.730 ;
        RECT  0.095 1.610 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  0.960 1.070 1.440 1.190 ;
        RECT  0.840 0.785 0.960 1.615 ;
        RECT  0.625 0.785 0.840 0.905 ;
        RECT  0.625 1.495 0.840 1.615 ;
        RECT  0.455 0.440 0.625 0.905 ;
        RECT  0.455 1.495 0.625 2.040 ;
    END
END BUFX8AD
MACRO CLKAND2X12AD
    CLASS CORE ;
    FOREIGN CLKAND2X12AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.370 0.670 3.565 2.065 ;
        RECT  3.340 0.805 3.370 2.065 ;
        RECT  2.805 0.805 3.340 1.615 ;
        RECT  2.635 0.670 2.805 2.065 ;
        RECT  2.525 0.805 2.635 1.615 ;
        RECT  2.085 0.805 2.525 0.935 ;
        RECT  2.100 1.375 2.525 1.615 ;
        RECT  1.915 1.375 2.100 2.090 ;
        RECT  1.915 0.670 2.085 0.935 ;
        END
        AntennaDiffArea 1.008 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.325 0.900 1.445 1.270 ;
        RECT  0.490 0.900 1.325 1.020 ;
        RECT  0.270 0.865 0.490 1.375 ;
        END
        AntennaGateArea 0.302 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.140 1.150 1.260 ;
        RECT  0.630 1.140 1.050 1.375 ;
        END
        AntennaGateArea 0.3029 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.950 -0.210 4.200 0.210 ;
        RECT  3.690 -0.210 3.950 0.710 ;
        RECT  3.210 -0.210 3.690 0.210 ;
        RECT  2.950 -0.210 3.210 0.685 ;
        RECT  2.490 -0.210 2.950 0.210 ;
        RECT  2.230 -0.210 2.490 0.685 ;
        RECT  1.660 -0.210 2.230 0.210 ;
        RECT  1.400 -0.210 1.660 0.540 ;
        RECT  0.380 -0.210 1.400 0.210 ;
        RECT  0.160 -0.210 0.380 0.720 ;
        RECT  0.000 -0.210 0.160 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.910 2.310 4.200 2.730 ;
        RECT  3.730 1.585 3.910 2.730 ;
        RECT  3.190 2.310 3.730 2.730 ;
        RECT  2.970 1.845 3.190 2.730 ;
        RECT  2.470 2.310 2.970 2.730 ;
        RECT  2.250 1.840 2.470 2.730 ;
        RECT  1.725 2.310 2.250 2.730 ;
        RECT  1.555 1.735 1.725 2.730 ;
        RECT  1.005 2.310 1.555 2.730 ;
        RECT  0.835 1.735 1.005 2.730 ;
        RECT  0.285 2.310 0.835 2.730 ;
        RECT  0.115 1.500 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  1.760 1.055 2.370 1.225 ;
        RECT  1.640 0.660 1.760 1.615 ;
        RECT  0.985 0.660 1.640 0.780 ;
        RECT  1.365 1.495 1.640 1.615 ;
        RECT  1.195 1.495 1.365 2.185 ;
        RECT  0.645 1.495 1.195 1.615 ;
        RECT  0.815 0.350 0.985 0.780 ;
        RECT  0.475 1.495 0.645 2.185 ;
    END
END CLKAND2X12AD
MACRO CLKAND2X2AD
    CLASS CORE ;
    FOREIGN CLKAND2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.625 1.330 2.165 ;
        RECT  1.135 0.625 1.190 0.795 ;
        RECT  1.160 1.385 1.190 2.165 ;
        END
        AntennaDiffArea 0.29 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.750 0.650 2.135 ;
        RECT  0.305 1.750 0.490 1.890 ;
        END
        AntennaGateArea 0.0577 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.240 1.280 ;
        RECT  0.070 1.020 0.210 1.650 ;
        END
        AntennaGateArea 0.0574 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.925 -0.210 1.400 0.210 ;
        RECT  0.705 -0.210 0.925 0.825 ;
        RECT  0.000 -0.210 0.705 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 2.310 1.400 2.730 ;
        RECT  0.775 1.455 0.945 2.730 ;
        RECT  0.370 2.310 0.775 2.730 ;
        RECT  0.110 2.040 0.370 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.555 1.010 0.980 1.270 ;
        RECT  0.385 0.675 0.555 1.585 ;
        RECT  0.090 0.675 0.385 0.845 ;
    END
END CLKAND2X2AD
MACRO CLKAND2X3AD
    CLASS CORE ;
    FOREIGN CLKAND2X3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.210 0.445 1.330 1.935 ;
        RECT  1.065 0.445 1.210 0.615 ;
        RECT  1.050 1.425 1.210 1.935 ;
        END
        AntennaDiffArea 0.295 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.020 0.810 1.375 ;
        END
        AntennaGateArea 0.0844 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.990 0.240 1.655 ;
        END
        AntennaGateArea 0.0844 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.910 -0.210 1.680 0.210 ;
        RECT  0.650 -0.210 0.910 0.615 ;
        RECT  0.000 -0.210 0.650 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.610 2.310 1.680 2.730 ;
        RECT  1.450 1.440 1.610 2.730 ;
        RECT  0.870 2.310 1.450 2.730 ;
        RECT  0.685 2.200 0.870 2.730 ;
        RECT  0.515 2.310 0.685 2.730 ;
        RECT  0.085 2.200 0.515 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  0.970 0.780 1.090 1.300 ;
        RECT  0.480 0.780 0.970 0.900 ;
        RECT  0.480 1.465 0.545 1.895 ;
        RECT  0.360 0.520 0.480 1.895 ;
        RECT  0.085 0.520 0.360 0.720 ;
    END
END CLKAND2X3AD
MACRO CLKAND2X4AD
    CLASS CORE ;
    FOREIGN CLKAND2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.325 0.550 1.450 2.165 ;
        RECT  1.195 0.550 1.325 0.745 ;
        RECT  1.190 1.285 1.325 2.165 ;
        END
        AntennaDiffArea 0.35 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 1.040 0.770 1.375 ;
        END
        AntennaGateArea 0.1123 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.045 0.410 1.205 ;
        RECT  0.070 1.045 0.210 1.375 ;
        END
        AntennaGateArea 0.112 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.745 -0.210 1.960 0.210 ;
        RECT  1.580 -0.210 1.745 0.790 ;
        RECT  0.990 -0.210 1.580 0.210 ;
        RECT  0.730 -0.210 0.990 0.660 ;
        RECT  0.000 -0.210 0.730 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.815 2.310 1.960 2.730 ;
        RECT  1.645 1.510 1.815 2.730 ;
        RECT  1.050 2.310 1.645 2.730 ;
        RECT  0.905 1.785 1.050 2.730 ;
        RECT  0.295 2.310 0.905 2.730 ;
        RECT  0.125 1.525 0.295 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.070 0.900 1.180 1.160 ;
        RECT  0.950 0.780 1.070 1.615 ;
        RECT  0.310 0.780 0.950 0.900 ;
        RECT  0.655 1.495 0.950 1.615 ;
        RECT  0.485 1.495 0.655 1.955 ;
        RECT  0.125 0.630 0.310 0.900 ;
    END
END CLKAND2X4AD
MACRO CLKAND2X6AD
    CLASS CORE ;
    FOREIGN CLKAND2X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.915 0.455 2.085 2.135 ;
        RECT  1.335 0.615 1.915 0.795 ;
        RECT  1.345 1.430 1.915 1.610 ;
        RECT  1.165 1.430 1.345 2.185 ;
        RECT  1.145 0.405 1.335 0.795 ;
        END
        AntennaDiffArea 0.618 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.805 1.375 ;
        END
        AntennaGateArea 0.151 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.240 1.375 ;
        END
        AntennaGateArea 0.151 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.750 -0.210 2.240 0.210 ;
        RECT  1.490 -0.210 1.750 0.495 ;
        RECT  0.970 -0.210 1.490 0.210 ;
        RECT  0.710 -0.210 0.970 0.730 ;
        RECT  0.000 -0.210 0.710 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.705 2.310 2.240 2.730 ;
        RECT  1.525 1.790 1.705 2.730 ;
        RECT  0.980 2.310 1.525 2.730 ;
        RECT  0.800 1.765 0.980 2.730 ;
        RECT  0.230 2.310 0.800 2.730 ;
        RECT  0.070 1.540 0.230 2.730 ;
        RECT  0.000 2.310 0.070 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.045 1.005 1.735 1.175 ;
        RECT  0.925 1.005 1.045 1.615 ;
        RECT  0.615 1.495 0.925 1.615 ;
        RECT  0.480 1.495 0.615 1.995 ;
        RECT  0.360 0.350 0.480 1.995 ;
        RECT  0.100 0.350 0.360 0.730 ;
    END
END CLKAND2X6AD
MACRO CLKAND2X8AD
    CLASS CORE ;
    FOREIGN CLKAND2X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.985 3.195 1.725 ;
        RECT  2.810 0.600 2.840 1.725 ;
        RECT  2.640 0.600 2.810 2.130 ;
        RECT  2.090 0.825 2.640 1.005 ;
        RECT  2.075 1.440 2.640 1.725 ;
        RECT  1.910 0.635 2.090 1.005 ;
        RECT  1.905 1.440 2.075 2.130 ;
        END
        AntennaDiffArea 0.668 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.315 0.900 1.435 1.270 ;
        RECT  0.440 0.900 1.315 1.020 ;
        RECT  0.210 0.900 0.440 1.070 ;
        RECT  0.070 0.855 0.210 1.375 ;
        END
        AntennaGateArea 0.218 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.140 1.140 1.375 ;
        END
        AntennaGateArea 0.2187 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.215 -0.210 3.360 0.210 ;
        RECT  2.965 -0.210 3.215 0.685 ;
        RECT  2.490 -0.210 2.965 0.210 ;
        RECT  2.230 -0.210 2.490 0.685 ;
        RECT  1.690 -0.210 2.230 0.210 ;
        RECT  1.430 -0.210 1.690 0.510 ;
        RECT  0.390 -0.210 1.430 0.210 ;
        RECT  0.130 -0.210 0.390 0.675 ;
        RECT  0.000 -0.210 0.130 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.175 2.310 3.360 2.730 ;
        RECT  2.995 1.845 3.175 2.730 ;
        RECT  2.445 2.310 2.995 2.730 ;
        RECT  2.275 1.845 2.445 2.730 ;
        RECT  1.740 2.310 2.275 2.730 ;
        RECT  1.520 1.750 1.740 2.730 ;
        RECT  1.020 2.310 1.520 2.730 ;
        RECT  0.800 1.750 1.020 2.730 ;
        RECT  0.280 2.310 0.800 2.730 ;
        RECT  0.100 1.520 0.280 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  1.750 1.140 2.520 1.260 ;
        RECT  1.630 0.630 1.750 1.615 ;
        RECT  0.975 0.630 1.630 0.750 ;
        RECT  1.355 1.495 1.630 1.615 ;
        RECT  1.185 1.495 1.355 1.950 ;
        RECT  0.650 1.495 1.185 1.615 ;
        RECT  0.805 0.505 0.975 0.750 ;
        RECT  0.530 1.495 0.650 1.950 ;
        RECT  0.465 1.520 0.530 1.950 ;
    END
END CLKAND2X8AD
MACRO CLKBUFX12AD
    CLASS CORE ;
    FOREIGN CLKBUFX12AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.595 0.685 2.795 2.070 ;
        RECT  2.075 0.685 2.595 1.675 ;
        RECT  1.905 0.445 2.075 2.070 ;
        RECT  1.885 0.685 1.905 1.660 ;
        RECT  1.355 0.685 1.885 0.885 ;
        RECT  1.385 1.375 1.885 1.660 ;
        RECT  1.185 1.375 1.385 2.065 ;
        RECT  1.185 0.415 1.355 0.885 ;
        END
        AntennaDiffArea 0.982 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.750 0.230 1.375 ;
        END
        AntennaGateArea 0.238 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.480 -0.210 3.360 0.210 ;
        RECT  2.220 -0.210 2.480 0.560 ;
        RECT  1.760 -0.210 2.220 0.210 ;
        RECT  1.500 -0.210 1.760 0.560 ;
        RECT  1.000 -0.210 1.500 0.210 ;
        RECT  0.820 -0.210 1.000 0.870 ;
        RECT  0.000 -0.210 0.820 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.155 2.310 3.360 2.730 ;
        RECT  2.985 1.585 3.155 2.730 ;
        RECT  2.435 2.310 2.985 2.730 ;
        RECT  2.265 1.845 2.435 2.730 ;
        RECT  1.715 2.310 2.265 2.730 ;
        RECT  1.545 1.845 1.715 2.730 ;
        RECT  0.995 2.310 1.545 2.730 ;
        RECT  0.825 1.495 0.995 2.730 ;
        RECT  0.275 2.310 0.825 2.730 ;
        RECT  0.105 1.495 0.275 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  0.635 1.075 1.705 1.195 ;
        RECT  0.515 0.445 0.635 2.100 ;
        RECT  0.465 0.445 0.515 0.875 ;
        RECT  0.465 1.410 0.515 2.100 ;
    END
END CLKBUFX12AD
MACRO CLKBUFX16AD
    CLASS CORE ;
    FOREIGN CLKBUFX16AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.650 0.815 3.810 2.120 ;
        RECT  3.265 0.815 3.650 1.630 ;
        RECT  3.115 0.505 3.265 1.630 ;
        RECT  3.095 0.505 3.115 2.075 ;
        RECT  2.945 0.575 3.095 2.075 ;
        RECT  2.545 0.575 2.945 1.630 ;
        RECT  2.395 0.505 2.545 1.630 ;
        RECT  2.375 0.505 2.395 2.065 ;
        RECT  2.290 0.575 2.375 2.065 ;
        RECT  1.825 0.575 2.290 0.775 ;
        RECT  2.225 1.245 2.290 2.065 ;
        RECT  1.675 1.245 2.225 1.630 ;
        RECT  1.655 0.505 1.825 0.775 ;
        RECT  1.505 1.245 1.675 2.065 ;
        END
        AntennaDiffArea 1.406 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 0.830 0.780 1.095 ;
        END
        AntennaGateArea 0.3168 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.630 -0.210 3.920 0.210 ;
        RECT  3.450 -0.210 3.630 0.525 ;
        RECT  2.910 -0.210 3.450 0.210 ;
        RECT  2.730 -0.210 2.910 0.445 ;
        RECT  2.190 -0.210 2.730 0.210 ;
        RECT  2.010 -0.210 2.190 0.445 ;
        RECT  1.390 -0.210 2.010 0.210 ;
        RECT  1.210 -0.210 1.390 0.675 ;
        RECT  0.595 -0.210 1.210 0.210 ;
        RECT  0.425 -0.210 0.595 0.565 ;
        RECT  0.000 -0.210 0.425 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.475 2.310 3.920 2.730 ;
        RECT  3.305 1.845 3.475 2.730 ;
        RECT  2.755 2.310 3.305 2.730 ;
        RECT  2.585 1.845 2.755 2.730 ;
        RECT  2.035 2.310 2.585 2.730 ;
        RECT  1.865 1.845 2.035 2.730 ;
        RECT  1.315 2.310 1.865 2.730 ;
        RECT  1.145 1.375 1.315 2.730 ;
        RECT  0.680 2.310 1.145 2.730 ;
        RECT  0.420 2.250 0.680 2.730 ;
        RECT  0.000 2.310 0.420 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  1.020 0.895 2.075 1.065 ;
        RECT  0.900 0.395 1.020 1.815 ;
        RECT  0.785 0.395 0.900 0.565 ;
        RECT  0.785 1.375 0.900 1.815 ;
        RECT  0.255 1.375 0.785 1.555 ;
        RECT  0.085 1.375 0.255 1.815 ;
    END
END CLKBUFX16AD
MACRO CLKBUFX1AD
    CLASS CORE ;
    FOREIGN CLKBUFX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.630 1.050 1.580 ;
        RECT  0.910 0.630 0.950 1.910 ;
        RECT  0.815 0.630 0.910 0.800 ;
        RECT  0.830 1.390 0.910 1.910 ;
        END
        AntennaDiffArea 0.179 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.145 0.420 1.280 ;
        RECT  0.070 1.145 0.210 1.375 ;
        END
        AntennaGateArea 0.0776 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.670 -0.210 1.120 0.210 ;
        RECT  0.410 -0.210 0.670 0.775 ;
        RECT  0.000 -0.210 0.410 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.640 2.310 1.120 2.730 ;
        RECT  0.420 1.765 0.640 2.730 ;
        RECT  0.000 2.310 0.420 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
        LAYER M1 ;
        RECT  0.570 0.895 0.690 1.625 ;
        RECT  0.265 0.895 0.570 1.015 ;
        RECT  0.255 1.505 0.570 1.625 ;
        RECT  0.095 0.585 0.265 1.015 ;
        RECT  0.085 1.505 0.255 1.935 ;
    END
END CLKBUFX1AD
MACRO CLKBUFX20AD
    CLASS CORE ;
    FOREIGN CLKBUFX20AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.405 0.890 4.575 2.065 ;
        RECT  3.855 0.890 4.405 1.725 ;
        RECT  3.685 0.505 3.855 2.085 ;
        RECT  3.135 0.890 3.685 1.725 ;
        RECT  3.135 0.460 3.180 0.720 ;
        RECT  2.965 0.460 3.135 2.080 ;
        RECT  2.920 0.460 2.965 1.725 ;
        RECT  2.525 0.585 2.920 1.725 ;
        RECT  2.415 0.585 2.525 0.890 ;
        RECT  2.415 1.385 2.525 1.725 ;
        RECT  2.245 0.505 2.415 0.890 ;
        RECT  2.245 1.385 2.415 2.075 ;
        RECT  1.695 0.585 2.245 0.890 ;
        RECT  1.695 1.385 2.245 1.725 ;
        RECT  1.525 0.505 1.695 0.890 ;
        RECT  1.525 1.385 1.695 2.075 ;
        END
        AntennaDiffArea 1.634 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 0.945 0.760 1.115 ;
        RECT  0.070 0.575 0.240 1.115 ;
        END
        AntennaGateArea 0.396 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.225 -0.210 5.040 0.210 ;
        RECT  4.045 -0.210 4.225 0.470 ;
        RECT  3.505 -0.210 4.045 0.210 ;
        RECT  3.325 -0.210 3.505 0.470 ;
        RECT  2.780 -0.210 3.325 0.210 ;
        RECT  2.600 -0.210 2.780 0.465 ;
        RECT  2.060 -0.210 2.600 0.210 ;
        RECT  1.880 -0.210 2.060 0.465 ;
        RECT  1.300 -0.210 1.880 0.210 ;
        RECT  1.120 -0.210 1.300 0.720 ;
        RECT  0.545 -0.210 1.120 0.210 ;
        RECT  0.375 -0.210 0.545 0.675 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.935 2.310 5.040 2.730 ;
        RECT  4.765 1.390 4.935 2.730 ;
        RECT  4.215 2.310 4.765 2.730 ;
        RECT  4.045 1.845 4.215 2.730 ;
        RECT  3.495 2.310 4.045 2.730 ;
        RECT  3.325 1.845 3.495 2.730 ;
        RECT  2.775 2.310 3.325 2.730 ;
        RECT  2.605 1.845 2.775 2.730 ;
        RECT  2.055 2.310 2.605 2.730 ;
        RECT  1.885 1.845 2.055 2.730 ;
        RECT  1.340 2.310 1.885 2.730 ;
        RECT  1.160 1.585 1.340 2.730 ;
        RECT  0.620 2.310 1.160 2.730 ;
        RECT  0.440 1.575 0.620 2.730 ;
        RECT  0.000 2.310 0.440 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.040 2.520 ;
        LAYER M1 ;
        RECT  1.000 1.085 2.340 1.205 ;
        RECT  0.950 0.630 1.000 2.065 ;
        RECT  0.880 0.330 0.950 2.065 ;
        RECT  0.690 0.330 0.880 0.750 ;
        RECT  0.805 1.315 0.880 2.065 ;
        RECT  0.255 1.315 0.805 1.435 ;
        RECT  0.085 1.315 0.255 2.095 ;
    END
END CLKBUFX20AD
MACRO CLKBUFX24AD
    CLASS CORE ;
    FOREIGN CLKBUFX24AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.995 0.390 5.040 0.650 ;
        RECT  4.825 0.390 4.995 2.125 ;
        RECT  4.780 0.390 4.825 1.445 ;
        RECT  4.275 0.540 4.780 1.445 ;
        RECT  4.105 0.435 4.275 2.140 ;
        RECT  3.555 0.540 4.105 1.445 ;
        RECT  3.385 0.435 3.555 2.150 ;
        RECT  2.955 0.540 3.385 1.445 ;
        RECT  2.835 0.540 2.955 0.720 ;
        RECT  2.835 1.195 2.955 1.445 ;
        RECT  2.665 0.435 2.835 0.720 ;
        RECT  2.665 1.195 2.835 2.145 ;
        RECT  2.120 0.540 2.665 0.720 ;
        RECT  2.115 1.195 2.665 1.445 ;
        RECT  1.940 0.355 2.120 0.720 ;
        RECT  1.945 1.195 2.115 2.070 ;
        END
        AntennaDiffArea 1.976 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.265 0.910 0.955 1.195 ;
        END
        AntennaGateArea 0.476 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.360 -0.210 5.600 0.210 ;
        RECT  5.180 -0.210 5.360 0.415 ;
        RECT  4.640 -0.210 5.180 0.210 ;
        RECT  4.460 -0.210 4.640 0.415 ;
        RECT  3.920 -0.210 4.460 0.210 ;
        RECT  3.740 -0.210 3.920 0.415 ;
        RECT  3.200 -0.210 3.740 0.210 ;
        RECT  3.020 -0.210 3.200 0.415 ;
        RECT  2.480 -0.210 3.020 0.210 ;
        RECT  2.300 -0.210 2.480 0.415 ;
        RECT  1.520 -0.210 2.300 0.210 ;
        RECT  1.340 -0.210 1.520 0.675 ;
        RECT  0.795 -0.210 1.340 0.210 ;
        RECT  0.615 -0.210 0.795 0.745 ;
        RECT  0.000 -0.210 0.615 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.355 2.310 5.600 2.730 ;
        RECT  5.185 1.585 5.355 2.730 ;
        RECT  4.635 2.310 5.185 2.730 ;
        RECT  4.465 1.585 4.635 2.730 ;
        RECT  3.915 2.310 4.465 2.730 ;
        RECT  3.745 1.585 3.915 2.730 ;
        RECT  3.195 2.310 3.745 2.730 ;
        RECT  3.025 1.585 3.195 2.730 ;
        RECT  2.475 2.310 3.025 2.730 ;
        RECT  2.305 1.585 2.475 2.730 ;
        RECT  1.760 2.310 2.305 2.730 ;
        RECT  1.580 1.465 1.760 2.730 ;
        RECT  1.040 2.310 1.580 2.730 ;
        RECT  0.860 1.735 1.040 2.730 ;
        RECT  0.320 2.310 0.860 2.730 ;
        RECT  0.140 1.415 0.320 2.730 ;
        RECT  0.000 2.310 0.140 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  1.220 0.840 2.775 1.010 ;
        RECT  1.225 1.360 1.395 2.065 ;
        RECT  1.220 1.360 1.225 1.540 ;
        RECT  1.150 0.655 1.220 1.540 ;
        RECT  1.100 0.345 1.150 1.540 ;
        RECT  0.980 0.345 1.100 0.775 ;
        RECT  0.675 1.360 1.100 1.540 ;
        RECT  0.505 1.360 0.675 2.190 ;
    END
END CLKBUFX24AD
MACRO CLKBUFX2AD
    CLASS CORE ;
    FOREIGN CLKBUFX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.535 1.050 2.140 ;
        RECT  0.855 0.535 0.910 0.705 ;
        RECT  0.880 1.360 0.910 2.140 ;
        END
        AntennaDiffArea 0.29 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.040 0.490 1.650 ;
        RECT  0.320 1.040 0.350 1.300 ;
        END
        AntennaGateArea 0.0777 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.710 -0.210 1.120 0.210 ;
        RECT  0.450 -0.210 0.710 0.680 ;
        RECT  0.000 -0.210 0.450 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.665 2.310 1.120 2.730 ;
        RECT  0.495 1.775 0.665 2.730 ;
        RECT  0.000 2.310 0.495 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
        LAYER M1 ;
        RECT  0.635 0.800 0.755 1.260 ;
        RECT  0.255 0.800 0.635 0.920 ;
        RECT  0.200 0.665 0.255 0.920 ;
        RECT  0.200 1.440 0.230 1.960 ;
        RECT  0.080 0.665 0.200 1.960 ;
    END
END CLKBUFX2AD
MACRO CLKBUFX32AD
    CLASS CORE ;
    FOREIGN CLKBUFX32AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.615 0.390 6.660 0.650 ;
        RECT  6.445 0.390 6.615 2.155 ;
        RECT  6.400 0.390 6.445 1.400 ;
        RECT  5.875 0.540 6.400 1.400 ;
        RECT  5.705 0.435 5.875 2.155 ;
        RECT  5.200 0.540 5.705 1.400 ;
        RECT  5.155 0.390 5.200 1.400 ;
        RECT  4.985 0.390 5.155 2.105 ;
        RECT  4.940 0.390 4.985 0.650 ;
        RECT  4.435 0.770 4.985 1.750 ;
        RECT  4.435 0.390 4.480 0.650 ;
        RECT  4.265 0.390 4.435 2.100 ;
        RECT  4.220 0.390 4.265 1.750 ;
        RECT  3.715 0.540 4.220 1.750 ;
        RECT  3.545 0.445 3.715 2.100 ;
        RECT  3.115 0.540 3.545 1.400 ;
        RECT  2.995 0.540 3.115 0.720 ;
        RECT  2.995 1.150 3.115 1.400 ;
        RECT  2.825 0.435 2.995 0.720 ;
        RECT  2.825 1.150 2.995 2.100 ;
        RECT  2.280 0.540 2.825 0.720 ;
        RECT  2.275 1.150 2.825 1.400 ;
        RECT  2.100 0.355 2.280 0.720 ;
        RECT  2.105 1.150 2.275 2.070 ;
        END
        AntennaDiffArea 2.745 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 0.795 1.235 0.965 ;
        RECT  0.545 0.795 1.115 1.095 ;
        END
        AntennaGateArea 0.62 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.240 -0.210 6.720 0.210 ;
        RECT  6.060 -0.210 6.240 0.415 ;
        RECT  5.520 -0.210 6.060 0.210 ;
        RECT  5.340 -0.210 5.520 0.415 ;
        RECT  4.800 -0.210 5.340 0.210 ;
        RECT  4.620 -0.210 4.800 0.415 ;
        RECT  4.080 -0.210 4.620 0.210 ;
        RECT  3.900 -0.210 4.080 0.415 ;
        RECT  3.360 -0.210 3.900 0.210 ;
        RECT  3.180 -0.210 3.360 0.415 ;
        RECT  2.640 -0.210 3.180 0.210 ;
        RECT  2.460 -0.210 2.640 0.415 ;
        RECT  1.925 -0.210 2.460 0.210 ;
        RECT  1.745 -0.210 1.925 0.415 ;
        RECT  1.200 -0.210 1.745 0.210 ;
        RECT  1.020 -0.210 1.200 0.420 ;
        RECT  0.480 -0.210 1.020 0.210 ;
        RECT  0.300 -0.210 0.480 0.420 ;
        RECT  0.000 -0.210 0.300 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.235 2.310 6.720 2.730 ;
        RECT  6.065 1.585 6.235 2.730 ;
        RECT  5.515 2.310 6.065 2.730 ;
        RECT  5.345 1.585 5.515 2.730 ;
        RECT  4.840 2.310 5.345 2.730 ;
        RECT  4.580 1.870 4.840 2.730 ;
        RECT  4.120 2.310 4.580 2.730 ;
        RECT  3.860 1.870 4.120 2.730 ;
        RECT  3.355 2.310 3.860 2.730 ;
        RECT  3.185 1.585 3.355 2.730 ;
        RECT  2.635 2.310 3.185 2.730 ;
        RECT  2.465 1.585 2.635 2.730 ;
        RECT  1.915 2.310 2.465 2.730 ;
        RECT  1.745 1.325 1.915 2.730 ;
        RECT  1.200 2.310 1.745 2.730 ;
        RECT  1.020 1.735 1.200 2.730 ;
        RECT  0.480 2.310 1.020 2.730 ;
        RECT  0.300 1.580 0.480 2.730 ;
        RECT  0.000 2.310 0.300 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.720 2.520 ;
        LAYER M1 ;
        RECT  1.555 0.840 2.980 0.960 ;
        RECT  1.435 0.455 1.555 2.065 ;
        RECT  1.385 0.455 1.435 0.670 ;
        RECT  1.385 1.360 1.435 2.065 ;
        RECT  0.835 0.550 1.385 0.670 ;
        RECT  0.835 1.360 1.385 1.540 ;
        RECT  0.665 0.455 0.835 0.670 ;
        RECT  0.665 1.360 0.835 2.190 ;
        RECT  0.620 0.550 0.665 0.670 ;
    END
END CLKBUFX32AD
MACRO CLKBUFX3AD
    CLASS CORE ;
    FOREIGN CLKBUFX3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.610 1.050 1.940 ;
        RECT  0.810 0.610 0.910 0.870 ;
        RECT  0.810 1.420 0.910 1.940 ;
        END
        AntennaDiffArea 0.246 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.065 0.420 1.235 ;
        RECT  0.070 1.065 0.210 1.375 ;
        END
        AntennaGateArea 0.0774 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.320 -0.210 1.400 0.210 ;
        RECT  1.170 -0.210 1.320 0.870 ;
        RECT  0.620 -0.210 1.170 0.210 ;
        RECT  0.360 -0.210 0.620 0.435 ;
        RECT  0.000 -0.210 0.360 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 2.310 1.400 2.730 ;
        RECT  1.290 1.470 1.330 2.730 ;
        RECT  1.170 1.450 1.290 2.730 ;
        RECT  0.620 2.310 1.170 2.730 ;
        RECT  0.360 2.200 0.620 2.730 ;
        RECT  0.000 2.310 0.360 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.690 1.030 0.780 1.290 ;
        RECT  0.570 0.705 0.690 1.685 ;
        RECT  0.085 0.705 0.570 0.875 ;
        RECT  0.085 1.515 0.570 1.685 ;
    END
END CLKBUFX3AD
MACRO CLKBUFX40AD
    CLASS CORE ;
    FOREIGN CLKBUFX40AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.575 0.380 7.620 0.640 ;
        RECT  7.405 0.380 7.575 2.165 ;
        RECT  7.360 0.380 7.405 1.400 ;
        RECT  6.855 0.540 7.360 1.400 ;
        RECT  6.685 0.435 6.855 2.095 ;
        RECT  6.135 0.540 6.685 1.400 ;
        RECT  5.965 0.435 6.135 2.105 ;
        RECT  5.460 0.540 5.965 1.400 ;
        RECT  5.415 0.390 5.460 1.400 ;
        RECT  5.245 0.390 5.415 2.100 ;
        RECT  5.200 0.390 5.245 0.650 ;
        RECT  4.695 0.770 5.245 1.750 ;
        RECT  4.525 0.455 4.695 2.100 ;
        RECT  3.975 0.535 4.525 1.750 ;
        RECT  3.805 0.435 3.975 2.100 ;
        RECT  3.255 0.535 3.805 0.705 ;
        RECT  3.255 1.150 3.805 1.400 ;
        RECT  3.085 0.435 3.255 0.705 ;
        RECT  3.085 1.150 3.255 2.100 ;
        RECT  2.535 0.535 3.085 0.705 ;
        RECT  2.535 1.150 3.085 1.400 ;
        RECT  2.365 0.355 2.535 0.705 ;
        RECT  2.365 1.150 2.535 2.100 ;
        END
        AntennaDiffArea 3.283 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.845 1.525 0.965 ;
        RECT  0.630 0.845 1.050 1.095 ;
        RECT  0.485 0.845 0.630 0.965 ;
        END
        AntennaGateArea 0.782 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.955 -0.210 8.120 0.210 ;
        RECT  7.785 -0.210 7.955 0.415 ;
        RECT  7.220 -0.210 7.785 0.210 ;
        RECT  7.040 -0.210 7.220 0.415 ;
        RECT  6.500 -0.210 7.040 0.210 ;
        RECT  6.320 -0.210 6.500 0.415 ;
        RECT  5.780 -0.210 6.320 0.210 ;
        RECT  5.600 -0.210 5.780 0.415 ;
        RECT  5.060 -0.210 5.600 0.210 ;
        RECT  4.880 -0.210 5.060 0.415 ;
        RECT  4.340 -0.210 4.880 0.210 ;
        RECT  4.160 -0.210 4.340 0.415 ;
        RECT  3.620 -0.210 4.160 0.210 ;
        RECT  3.440 -0.210 3.620 0.415 ;
        RECT  2.900 -0.210 3.440 0.210 ;
        RECT  2.720 -0.210 2.900 0.415 ;
        RECT  2.185 -0.210 2.720 0.210 ;
        RECT  2.005 -0.210 2.185 0.415 ;
        RECT  1.460 -0.210 2.005 0.210 ;
        RECT  1.280 -0.210 1.460 0.415 ;
        RECT  0.740 -0.210 1.280 0.210 ;
        RECT  0.560 -0.210 0.740 0.415 ;
        RECT  0.000 -0.210 0.560 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.955 2.310 8.120 2.730 ;
        RECT  7.785 1.465 7.955 2.730 ;
        RECT  7.215 2.310 7.785 2.730 ;
        RECT  7.045 1.585 7.215 2.730 ;
        RECT  6.495 2.310 7.045 2.730 ;
        RECT  6.325 1.585 6.495 2.730 ;
        RECT  5.775 2.310 6.325 2.730 ;
        RECT  5.605 1.585 5.775 2.730 ;
        RECT  5.100 2.310 5.605 2.730 ;
        RECT  4.840 1.870 5.100 2.730 ;
        RECT  4.380 2.310 4.840 2.730 ;
        RECT  4.120 1.870 4.380 2.730 ;
        RECT  3.615 2.310 4.120 2.730 ;
        RECT  3.445 1.585 3.615 2.730 ;
        RECT  2.895 2.310 3.445 2.730 ;
        RECT  2.725 1.585 2.895 2.730 ;
        RECT  2.175 2.310 2.725 2.730 ;
        RECT  2.005 1.325 2.175 2.730 ;
        RECT  1.460 2.310 2.005 2.730 ;
        RECT  1.280 1.735 1.460 2.730 ;
        RECT  0.740 2.310 1.280 2.730 ;
        RECT  0.560 1.735 0.740 2.730 ;
        RECT  0.000 2.310 0.560 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.120 2.520 ;
        LAYER M1 ;
        RECT  1.815 0.830 3.600 0.950 ;
        RECT  1.645 0.455 1.815 2.065 ;
        RECT  1.095 0.535 1.645 0.695 ;
        RECT  1.095 1.360 1.645 1.540 ;
        RECT  0.925 0.455 1.095 0.695 ;
        RECT  0.925 1.360 1.095 2.190 ;
        RECT  0.375 0.535 0.925 0.695 ;
        RECT  0.375 1.360 0.925 1.540 ;
        RECT  0.205 0.455 0.375 0.695 ;
        RECT  0.205 1.360 0.375 2.190 ;
    END
END CLKBUFX40AD
MACRO CLKBUFX4AD
    CLASS CORE ;
    FOREIGN CLKBUFX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.955 0.630 1.050 1.705 ;
        RECT  0.910 0.630 0.955 2.165 ;
        RECT  0.810 0.630 0.910 0.890 ;
        RECT  0.785 1.475 0.910 2.165 ;
        END
        AntennaDiffArea 0.328 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.070 0.400 1.235 ;
        RECT  0.070 1.070 0.210 1.375 ;
        END
        AntennaGateArea 0.0794 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 -0.210 1.400 0.210 ;
        RECT  1.170 -0.210 1.330 0.875 ;
        RECT  0.610 -0.210 1.170 0.210 ;
        RECT  0.350 -0.210 0.610 0.400 ;
        RECT  0.000 -0.210 0.350 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.330 2.310 1.400 2.730 ;
        RECT  1.170 1.435 1.330 2.730 ;
        RECT  0.570 2.310 1.170 2.730 ;
        RECT  0.540 2.230 0.570 2.730 ;
        RECT  0.320 2.200 0.540 2.730 ;
        RECT  0.310 2.230 0.320 2.730 ;
        RECT  0.000 2.310 0.310 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.665 1.030 0.780 1.290 ;
        RECT  0.545 0.755 0.665 1.615 ;
        RECT  0.255 0.755 0.545 0.875 ;
        RECT  0.255 1.495 0.545 1.615 ;
        RECT  0.085 0.705 0.255 0.875 ;
        RECT  0.085 1.495 0.255 1.925 ;
    END
END CLKBUFX4AD
MACRO CLKBUFX6AD
    CLASS CORE ;
    FOREIGN CLKBUFX6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.765 0.770 1.890 1.655 ;
        RECT  1.720 0.770 1.765 2.170 ;
        RECT  1.215 0.770 1.720 0.950 ;
        RECT  1.595 1.455 1.720 2.170 ;
        RECT  1.045 1.455 1.595 1.615 ;
        RECT  1.045 0.475 1.215 0.950 ;
        RECT  0.875 1.455 1.045 2.165 ;
        END
        AntennaDiffArea 0.594 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.090 0.515 1.250 ;
        RECT  0.070 1.090 0.210 1.375 ;
        END
        AntennaGateArea 0.119 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.630 -0.210 1.960 0.210 ;
        RECT  1.370 -0.210 1.630 0.650 ;
        RECT  0.890 -0.210 1.370 0.210 ;
        RECT  0.630 -0.210 0.890 0.650 ;
        RECT  0.000 -0.210 0.630 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.410 2.310 1.960 2.730 ;
        RECT  1.230 1.735 1.410 2.730 ;
        RECT  0.690 2.310 1.230 2.730 ;
        RECT  0.510 1.735 0.690 2.730 ;
        RECT  0.000 2.310 0.510 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.460 1.110 1.490 1.230 ;
        RECT  0.755 1.110 1.460 1.285 ;
        RECT  0.635 0.785 0.755 1.615 ;
        RECT  0.395 0.785 0.635 0.905 ;
        RECT  0.305 1.495 0.635 1.615 ;
        RECT  0.225 0.735 0.395 0.905 ;
        RECT  0.135 1.495 0.305 2.010 ;
    END
END CLKBUFX6AD
MACRO CLKBUFX8AD
    CLASS CORE ;
    FOREIGN CLKBUFX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.065 0.660 2.110 2.035 ;
        RECT  1.895 0.660 2.065 2.110 ;
        RECT  1.875 0.660 1.895 2.035 ;
        RECT  1.610 0.660 1.875 1.630 ;
        RECT  1.100 0.660 1.610 0.920 ;
        RECT  1.345 1.400 1.610 1.630 ;
        RECT  1.175 1.400 1.345 2.110 ;
        END
        AntennaDiffArea 0.709 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.065 0.730 1.235 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.1597 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.720 -0.210 2.520 0.210 ;
        RECT  1.460 -0.210 1.720 0.540 ;
        RECT  0.940 -0.210 1.460 0.210 ;
        RECT  0.680 -0.210 0.940 0.700 ;
        RECT  0.000 -0.210 0.680 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.425 2.310 2.520 2.730 ;
        RECT  2.255 1.585 2.425 2.730 ;
        RECT  1.705 2.310 2.255 2.730 ;
        RECT  1.535 1.750 1.705 2.730 ;
        RECT  0.985 2.310 1.535 2.730 ;
        RECT  0.815 1.680 0.985 2.730 ;
        RECT  0.330 2.310 0.815 2.730 ;
        RECT  0.130 2.205 0.330 2.730 ;
        RECT  0.000 2.310 0.130 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  0.970 1.110 1.450 1.230 ;
        RECT  0.850 0.825 0.970 1.530 ;
        RECT  0.530 0.825 0.850 0.945 ;
        RECT  0.595 1.400 0.850 1.530 ;
        RECT  0.425 1.400 0.595 1.830 ;
        RECT  0.330 0.680 0.530 0.945 ;
    END
END CLKBUFX8AD
MACRO CLKINVX12AD
    CLASS CORE ;
    FOREIGN CLKINVX12AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.015 0.890 2.055 2.090 ;
        RECT  1.885 0.465 2.015 2.090 ;
        RECT  1.845 0.465 1.885 1.630 ;
        RECT  1.335 0.890 1.845 1.630 ;
        RECT  1.295 0.890 1.335 2.090 ;
        RECT  1.165 0.465 1.295 2.090 ;
        RECT  1.125 0.465 1.165 1.630 ;
        RECT  0.615 1.400 1.125 1.630 ;
        RECT  0.445 1.400 0.615 2.090 ;
        RECT  0.440 1.400 0.445 1.630 ;
        END
        AntennaDiffArea 0.982 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.110 0.800 1.230 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.754 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.380 -0.210 2.520 0.210 ;
        RECT  2.200 -0.210 2.380 0.640 ;
        RECT  1.660 -0.210 2.200 0.210 ;
        RECT  1.480 -0.210 1.660 0.640 ;
        RECT  0.935 -0.210 1.480 0.210 ;
        RECT  0.765 -0.210 0.935 0.895 ;
        RECT  0.000 -0.210 0.765 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.415 2.310 2.520 2.730 ;
        RECT  2.245 1.660 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 1.760 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.760 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.560 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
	 END
END CLKINVX12AD
MACRO CLKINVX16AD
    CLASS CORE ;
    FOREIGN CLKINVX16AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.605 1.375 2.775 2.065 ;
        RECT  2.235 1.375 2.605 1.685 ;
        RECT  2.205 0.610 2.235 1.685 ;
        RECT  2.055 0.455 2.205 1.685 ;
        RECT  2.035 0.455 2.055 2.065 ;
        RECT  1.885 0.610 2.035 2.065 ;
        RECT  1.425 0.610 1.885 1.685 ;
        RECT  1.335 0.455 1.425 1.685 ;
        RECT  1.290 0.455 1.335 2.065 ;
        RECT  1.255 0.455 1.290 0.890 ;
        RECT  1.165 1.375 1.290 2.065 ;
        RECT  0.645 0.610 1.255 0.890 ;
        RECT  0.615 1.375 1.165 1.685 ;
        RECT  0.475 0.455 0.645 0.890 ;
        RECT  0.445 1.375 0.615 2.065 ;
        END
        AntennaDiffArea 1.36 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.060 1.080 1.200 ;
        RECT  0.070 0.585 0.210 1.200 ;
        END
        AntennaGateArea 1.006 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.570 -0.210 3.360 0.210 ;
        RECT  2.390 -0.210 2.570 0.885 ;
        RECT  1.860 -0.210 2.390 0.210 ;
        RECT  1.600 -0.210 1.860 0.490 ;
        RECT  1.080 -0.210 1.600 0.210 ;
        RECT  0.820 -0.210 1.080 0.490 ;
        RECT  0.000 -0.210 0.820 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.135 2.310 3.360 2.730 ;
        RECT  2.965 1.375 3.135 2.730 ;
        RECT  2.415 2.310 2.965 2.730 ;
        RECT  2.245 1.845 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 1.845 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.845 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.375 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
	 END
END CLKINVX16AD
MACRO CLKINVX1AD
    CLASS CORE ;
    FOREIGN CLKINVX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.725 0.585 0.770 1.095 ;
        RECT  0.685 0.585 0.725 1.625 ;
        RECT  0.605 0.575 0.685 1.925 ;
        RECT  0.515 0.575 0.605 0.745 ;
        RECT  0.515 1.495 0.605 1.925 ;
        END
        AntennaDiffArea 0.183 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.085 0.420 1.240 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.077 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.325 -0.210 0.840 0.210 ;
        RECT  0.155 -0.210 0.325 0.745 ;
        RECT  0.000 -0.210 0.155 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.325 2.310 0.840 2.730 ;
        RECT  0.155 1.495 0.325 2.730 ;
        RECT  0.000 2.310 0.155 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 0.840 2.520 ;
	 END
END CLKINVX1AD
MACRO CLKINVX20AD
    CLASS CORE ;
    FOREIGN CLKINVX20AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.360 0.510 3.520 2.110 ;
        RECT  3.095 0.510 3.360 1.430 ;
        RECT  2.925 0.375 3.095 1.430 ;
        RECT  2.775 0.510 2.925 1.430 ;
        RECT  2.605 0.510 2.775 2.065 ;
        RECT  2.355 0.510 2.605 1.430 ;
        RECT  2.185 0.375 2.355 1.430 ;
        RECT  2.055 0.510 2.185 1.430 ;
        RECT  1.885 0.510 2.055 2.065 ;
        RECT  1.625 0.510 1.885 1.685 ;
        RECT  1.455 0.375 1.625 1.685 ;
        RECT  1.335 0.510 1.455 1.685 ;
        RECT  1.285 0.510 1.335 2.065 ;
        RECT  0.885 0.510 1.285 0.690 ;
        RECT  1.165 1.375 1.285 2.065 ;
        RECT  0.615 1.375 1.165 1.685 ;
        RECT  0.715 0.375 0.885 0.690 ;
        RECT  0.445 1.375 0.615 2.065 ;
        END
        AntennaDiffArea 1.764 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.895 1.095 1.095 ;
        RECT  0.070 0.585 0.210 1.095 ;
        END
        AntennaGateArea 1.26 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.510 -0.210 3.640 0.210 ;
        RECT  3.250 -0.210 3.510 0.390 ;
        RECT  2.770 -0.210 3.250 0.210 ;
        RECT  2.510 -0.210 2.770 0.390 ;
        RECT  2.040 -0.210 2.510 0.210 ;
        RECT  1.780 -0.210 2.040 0.390 ;
        RECT  1.300 -0.210 1.780 0.210 ;
        RECT  1.040 -0.210 1.300 0.390 ;
        RECT  0.520 -0.210 1.040 0.210 ;
        RECT  0.340 -0.210 0.520 0.545 ;
        RECT  0.000 -0.210 0.340 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.135 2.310 3.640 2.730 ;
        RECT  2.965 1.585 3.135 2.730 ;
        RECT  2.415 2.310 2.965 2.730 ;
        RECT  2.245 1.585 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 1.845 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.845 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.375 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
	 END
END CLKINVX20AD
MACRO CLKINVX24AD
    CLASS CORE ;
    FOREIGN CLKINVX24AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.095 0.510 4.265 2.115 ;
        RECT  3.805 0.510 4.095 1.430 ;
        RECT  3.635 0.375 3.805 1.430 ;
        RECT  3.495 0.510 3.635 1.430 ;
        RECT  3.325 0.510 3.495 2.065 ;
        RECT  3.075 0.510 3.325 1.430 ;
        RECT  2.905 0.375 3.075 1.430 ;
        RECT  2.775 0.510 2.905 1.430 ;
        RECT  2.605 0.510 2.775 2.065 ;
        RECT  2.355 0.510 2.605 1.430 ;
        RECT  2.185 0.375 2.355 1.430 ;
        RECT  2.055 0.510 2.185 1.430 ;
        RECT  1.885 0.510 2.055 2.065 ;
        RECT  1.625 0.510 1.885 1.685 ;
        RECT  1.455 0.375 1.625 1.685 ;
        RECT  1.335 0.510 1.455 1.685 ;
        RECT  1.255 0.510 1.335 2.065 ;
        RECT  0.885 0.510 1.255 0.835 ;
        RECT  1.165 1.375 1.255 2.065 ;
        RECT  0.615 1.375 1.165 1.685 ;
        RECT  0.715 0.375 0.885 0.835 ;
        RECT  0.445 1.375 0.615 2.065 ;
        END
        AntennaDiffArea 2.076 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.005 1.095 1.175 ;
        RECT  0.070 0.585 0.210 1.175 ;
        END
        AntennaGateArea 1.5062 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.220 -0.210 4.480 0.210 ;
        RECT  3.960 -0.210 4.220 0.390 ;
        RECT  3.480 -0.210 3.960 0.210 ;
        RECT  3.220 -0.210 3.480 0.390 ;
        RECT  2.760 -0.210 3.220 0.210 ;
        RECT  2.500 -0.210 2.760 0.390 ;
        RECT  2.040 -0.210 2.500 0.210 ;
        RECT  1.780 -0.210 2.040 0.390 ;
        RECT  1.300 -0.210 1.780 0.210 ;
        RECT  1.040 -0.210 1.300 0.390 ;
        RECT  0.520 -0.210 1.040 0.210 ;
        RECT  0.340 -0.210 0.520 0.415 ;
        RECT  0.000 -0.210 0.340 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.855 2.310 4.480 2.730 ;
        RECT  3.685 1.585 3.855 2.730 ;
        RECT  3.135 2.310 3.685 2.730 ;
        RECT  2.965 1.585 3.135 2.730 ;
        RECT  2.415 2.310 2.965 2.730 ;
        RECT  2.245 1.585 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 1.845 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.845 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.375 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
	 END
END CLKINVX24AD
MACRO CLKINVX2AD
    CLASS CORE ;
    FOREIGN CLKINVX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.675 0.585 0.770 0.815 ;
        RECT  0.525 0.585 0.675 2.110 ;
        RECT  0.350 0.585 0.525 0.815 ;
        RECT  0.445 1.420 0.525 2.110 ;
        END
        AntennaDiffArea 0.29 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.050 0.400 1.210 ;
        RECT  0.070 1.050 0.210 1.655 ;
        END
        AntennaGateArea 0.126 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.230 -0.210 0.840 0.210 ;
        RECT  0.070 -0.210 0.230 0.880 ;
        RECT  0.000 -0.210 0.070 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.255 2.310 0.840 2.730 ;
        RECT  0.085 1.775 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 0.840 2.520 ;
	 END
END CLKINVX2AD
MACRO CLKINVX32AD
    CLASS CORE ;
    FOREIGN CLKINVX32AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.475 0.330 5.520 0.590 ;
        RECT  5.260 0.330 5.475 1.470 ;
        RECT  4.935 0.490 5.260 1.470 ;
        RECT  4.765 0.490 4.935 2.065 ;
        RECT  4.615 0.490 4.765 1.470 ;
        RECT  4.445 0.375 4.615 1.470 ;
        RECT  4.215 0.490 4.445 1.470 ;
        RECT  4.045 0.490 4.215 2.065 ;
        RECT  3.755 0.490 4.045 1.420 ;
        RECT  3.585 0.375 3.755 1.420 ;
        RECT  3.495 0.510 3.585 1.420 ;
        RECT  3.325 0.510 3.495 2.065 ;
        RECT  3.035 0.510 3.325 1.420 ;
        RECT  2.865 0.375 3.035 1.420 ;
        RECT  2.775 0.510 2.865 1.420 ;
        RECT  2.605 0.510 2.775 2.065 ;
        RECT  2.315 0.510 2.605 1.420 ;
        RECT  2.145 0.375 2.315 1.420 ;
        RECT  2.055 0.510 2.145 1.420 ;
        RECT  1.885 0.510 2.055 2.065 ;
        RECT  1.595 0.510 1.885 1.675 ;
        RECT  1.425 0.375 1.595 1.675 ;
        RECT  1.335 0.510 1.425 1.675 ;
        RECT  1.255 0.510 1.335 2.100 ;
        RECT  0.875 0.510 1.255 0.825 ;
        RECT  1.165 1.365 1.255 2.100 ;
        RECT  0.615 1.365 1.165 1.675 ;
        RECT  0.705 0.375 0.875 0.825 ;
        RECT  0.445 1.365 0.615 2.100 ;
        END
        AntennaDiffArea 2.729 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.005 1.095 1.175 ;
        RECT  0.070 0.585 0.210 1.175 ;
        END
        AntennaGateArea 2.0102 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.090 -0.210 5.600 0.210 ;
        RECT  4.830 -0.210 5.090 0.335 ;
        RECT  4.230 -0.210 4.830 0.210 ;
        RECT  3.970 -0.210 4.230 0.335 ;
        RECT  3.440 -0.210 3.970 0.210 ;
        RECT  3.180 -0.210 3.440 0.390 ;
        RECT  2.720 -0.210 3.180 0.210 ;
        RECT  2.460 -0.210 2.720 0.390 ;
        RECT  2.000 -0.210 2.460 0.210 ;
        RECT  1.740 -0.210 2.000 0.390 ;
        RECT  1.280 -0.210 1.740 0.210 ;
        RECT  1.020 -0.210 1.280 0.390 ;
        RECT  0.525 -0.210 1.020 0.210 ;
        RECT  0.345 -0.210 0.525 0.545 ;
        RECT  0.000 -0.210 0.345 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.345 2.310 5.600 2.730 ;
        RECT  5.175 1.670 5.345 2.730 ;
        RECT  4.575 2.310 5.175 2.730 ;
        RECT  4.405 1.845 4.575 2.730 ;
        RECT  3.855 2.310 4.405 2.730 ;
        RECT  3.685 1.585 3.855 2.730 ;
        RECT  3.135 2.310 3.685 2.730 ;
        RECT  2.965 1.585 3.135 2.730 ;
        RECT  2.415 2.310 2.965 2.730 ;
        RECT  2.245 1.845 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 1.845 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.845 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.410 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
	 END
END CLKINVX32AD
MACRO CLKINVX3AD
    CLASS CORE ;
    FOREIGN CLKINVX3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 0.635 0.770 1.100 ;
        RECT  0.505 0.635 0.680 1.865 ;
        RECT  0.475 1.435 0.505 1.865 ;
        END
        AntennaDiffArea 0.295 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.100 0.355 1.260 ;
        RECT  0.070 1.100 0.210 1.655 ;
        END
        AntennaGateArea 0.189 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.355 -0.210 1.120 0.210 ;
        RECT  0.185 -0.210 0.355 0.905 ;
        RECT  0.000 -0.210 0.185 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.010 2.310 1.120 2.730 ;
        RECT  0.835 1.455 1.010 2.730 ;
        RECT  0.285 2.310 0.835 2.730 ;
        RECT  0.115 1.775 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
	 END
END CLKINVX3AD
MACRO CLKINVX40AD
    CLASS CORE ;
    FOREIGN CLKINVX40AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.210 0.510 6.380 2.155 ;
        RECT  6.060 0.510 6.210 1.420 ;
        RECT  5.890 0.375 6.060 1.420 ;
        RECT  5.660 0.510 5.890 1.420 ;
        RECT  5.490 0.510 5.660 2.065 ;
        RECT  5.340 0.510 5.490 1.420 ;
        RECT  5.170 0.375 5.340 1.420 ;
        RECT  4.940 0.510 5.170 1.420 ;
        RECT  4.770 0.510 4.940 2.065 ;
        RECT  4.615 0.510 4.770 1.420 ;
        RECT  4.445 0.375 4.615 1.420 ;
        RECT  4.220 0.510 4.445 1.420 ;
        RECT  4.050 0.510 4.220 2.065 ;
        RECT  3.895 0.510 4.050 1.420 ;
        RECT  3.725 0.375 3.895 1.420 ;
        RECT  3.500 0.510 3.725 1.420 ;
        RECT  3.330 0.510 3.500 2.065 ;
        RECT  3.225 0.510 3.330 1.470 ;
        RECT  3.175 0.490 3.225 1.470 ;
        RECT  3.005 0.375 3.175 1.470 ;
        RECT  2.775 0.490 3.005 1.470 ;
        RECT  2.605 0.490 2.775 2.065 ;
        RECT  2.315 0.490 2.605 1.705 ;
        RECT  2.145 0.375 2.315 1.705 ;
        RECT  2.095 0.490 2.145 1.705 ;
        RECT  2.070 0.510 2.095 1.705 ;
        RECT  1.595 0.510 2.070 0.795 ;
        RECT  2.055 1.365 2.070 1.705 ;
        RECT  1.885 1.365 2.055 2.065 ;
        RECT  1.335 1.365 1.885 1.705 ;
        RECT  1.425 0.375 1.595 0.795 ;
        RECT  0.875 0.510 1.425 0.795 ;
        RECT  1.165 1.365 1.335 2.100 ;
        RECT  0.615 1.365 1.165 1.705 ;
        RECT  0.705 0.375 0.875 0.795 ;
        RECT  0.445 1.365 0.615 2.100 ;
        END
        AntennaDiffArea 3.268 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.970 1.890 1.115 ;
        RECT  0.070 0.605 0.210 1.115 ;
        END
        AntennaGateArea 2.513 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.465 -0.210 7.000 0.210 ;
        RECT  6.205 -0.210 6.465 0.390 ;
        RECT  5.745 -0.210 6.205 0.210 ;
        RECT  5.485 -0.210 5.745 0.390 ;
        RECT  5.025 -0.210 5.485 0.210 ;
        RECT  4.765 -0.210 5.025 0.390 ;
        RECT  4.300 -0.210 4.765 0.210 ;
        RECT  4.040 -0.210 4.300 0.390 ;
        RECT  3.580 -0.210 4.040 0.210 ;
        RECT  3.320 -0.210 3.580 0.390 ;
        RECT  2.790 -0.210 3.320 0.210 ;
        RECT  2.530 -0.210 2.790 0.350 ;
        RECT  2.000 -0.210 2.530 0.210 ;
        RECT  1.740 -0.210 2.000 0.390 ;
        RECT  1.280 -0.210 1.740 0.210 ;
        RECT  1.020 -0.210 1.280 0.390 ;
        RECT  0.525 -0.210 1.020 0.210 ;
        RECT  0.345 -0.210 0.525 0.545 ;
        RECT  0.000 -0.210 0.345 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.740 2.310 7.000 2.730 ;
        RECT  6.570 1.715 6.740 2.730 ;
        RECT  6.020 2.310 6.570 2.730 ;
        RECT  5.850 1.715 6.020 2.730 ;
        RECT  5.300 2.310 5.850 2.730 ;
        RECT  5.130 1.585 5.300 2.730 ;
        RECT  4.580 2.310 5.130 2.730 ;
        RECT  4.410 1.585 4.580 2.730 ;
        RECT  3.860 2.310 4.410 2.730 ;
        RECT  3.690 1.585 3.860 2.730 ;
        RECT  3.180 2.310 3.690 2.730 ;
        RECT  2.920 1.610 3.180 2.730 ;
        RECT  2.415 2.310 2.920 2.730 ;
        RECT  2.245 1.845 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 1.845 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.845 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.410 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
	 END
END CLKINVX40AD
MACRO CLKINVX4AD
    CLASS CORE ;
    FOREIGN CLKINVX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.645 1.005 0.770 1.515 ;
        RECT  0.515 0.690 0.645 2.120 ;
        RECT  0.475 0.690 0.515 0.860 ;
        RECT  0.475 1.430 0.515 2.120 ;
        END
        AntennaDiffArea 0.328 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.085 0.395 1.225 ;
        RECT  0.070 1.085 0.210 1.655 ;
        END
        AntennaGateArea 0.252 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 -0.210 1.120 0.210 ;
        RECT  0.890 -0.210 1.050 0.860 ;
        RECT  0.285 -0.210 0.890 0.210 ;
        RECT  0.115 -0.210 0.285 0.860 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.005 2.310 1.120 2.730 ;
        RECT  0.835 1.695 1.005 2.730 ;
        RECT  0.285 2.310 0.835 2.730 ;
        RECT  0.115 1.845 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
	 END
END CLKINVX4AD
MACRO CLKINVX6AD
    CLASS CORE ;
    FOREIGN CLKINVX6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.145 1.430 2.000 ;
        RECT  1.125 1.145 1.190 1.600 ;
        RECT  0.975 0.475 1.125 1.600 ;
        RECT  0.895 0.475 0.975 0.905 ;
        RECT  0.665 1.360 0.975 1.600 ;
        RECT  0.495 1.360 0.665 1.990 ;
        END
        AntennaDiffArea 0.584 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.110 0.850 1.230 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.377 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.465 -0.210 1.680 0.210 ;
        RECT  1.255 -0.210 1.465 0.875 ;
        RECT  0.705 -0.210 1.255 0.210 ;
        RECT  0.535 -0.210 0.705 0.900 ;
        RECT  0.000 -0.210 0.535 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.045 2.310 1.680 2.730 ;
        RECT  0.875 1.730 1.045 2.730 ;
        RECT  0.305 2.310 0.875 2.730 ;
        RECT  0.135 1.540 0.305 2.730 ;
        RECT  0.000 2.310 0.135 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
	 END
END CLKINVX6AD
MACRO CLKINVX8AD
    CLASS CORE ;
    FOREIGN CLKINVX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.760 1.545 0.880 ;
        RECT  1.385 0.740 1.470 1.515 ;
        RECT  1.195 0.740 1.385 1.955 ;
        RECT  0.980 0.740 1.195 1.595 ;
        RECT  0.655 0.740 0.980 0.905 ;
        RECT  0.670 1.350 0.980 1.595 ;
        RECT  0.470 1.350 0.670 2.085 ;
        RECT  0.485 0.475 0.655 0.905 ;
        END
        AntennaDiffArea 0.694 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.820 1.110 0.840 1.230 ;
        RECT  0.210 1.100 0.820 1.230 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.503 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.090 -0.210 1.960 0.210 ;
        RECT  0.830 -0.210 1.090 0.620 ;
        RECT  0.295 -0.210 0.830 0.210 ;
        RECT  0.125 -0.210 0.295 0.740 ;
        RECT  0.000 -0.210 0.125 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 2.310 1.960 2.730 ;
        RECT  1.590 1.540 1.765 2.730 ;
        RECT  1.015 2.310 1.590 2.730 ;
        RECT  0.845 1.735 1.015 2.730 ;
        RECT  0.295 2.310 0.845 2.730 ;
        RECT  0.125 1.555 0.295 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
	 END
END CLKINVX8AD
MACRO CLKMX2X12AD
    CLASS CORE ;
    FOREIGN CLKMX2X12AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.255 0.705 4.430 2.110 ;
        RECT  3.655 0.705 4.255 1.875 ;
        RECT  3.485 0.425 3.655 2.145 ;
        RECT  2.895 0.705 3.485 0.940 ;
        RECT  2.980 1.455 3.485 1.875 ;
        RECT  2.830 1.455 2.980 2.050 ;
        RECT  2.710 0.435 2.895 0.940 ;
        RECT  2.765 1.620 2.830 2.050 ;
        END
        AntennaDiffArea 1.038 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.465 0.990 1.585 1.870 ;
        RECT  0.240 1.750 1.465 1.870 ;
        RECT  0.240 2.070 0.345 2.190 ;
        RECT  0.070 1.705 0.240 2.190 ;
        END
        AntennaGateArea 0.193 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.820 1.150 ;
        END
        AntennaGateArea 0.126 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 0.865 2.450 1.260 ;
        END
        AntennaGateArea 0.126 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.070 -0.210 5.040 0.210 ;
        RECT  3.810 -0.210 4.070 0.570 ;
        RECT  3.340 -0.210 3.810 0.210 ;
        RECT  3.080 -0.210 3.340 0.570 ;
        RECT  2.560 -0.210 3.080 0.210 ;
        RECT  2.300 -0.210 2.560 0.730 ;
        RECT  0.645 -0.210 2.300 0.210 ;
        RECT  0.475 -0.210 0.645 0.495 ;
        RECT  0.000 -0.210 0.475 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.785 2.310 5.040 2.730 ;
        RECT  4.615 1.420 4.785 2.730 ;
        RECT  4.035 2.310 4.615 2.730 ;
        RECT  3.865 1.995 4.035 2.730 ;
        RECT  3.295 2.310 3.865 2.730 ;
        RECT  3.125 1.995 3.295 2.730 ;
        RECT  2.600 2.310 3.125 2.730 ;
        RECT  2.430 1.800 2.600 2.730 ;
        RECT  0.655 2.310 2.430 2.730 ;
        RECT  0.485 1.990 0.655 2.730 ;
        RECT  0.000 2.310 0.485 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.040 2.520 ;
        LAYER M1 ;
        RECT  2.705 1.115 3.365 1.235 ;
        RECT  2.585 1.115 2.705 1.500 ;
        RECT  2.310 1.380 2.585 1.500 ;
        RECT  2.190 1.380 2.310 2.140 ;
        RECT  1.825 2.020 2.190 2.140 ;
        RECT  1.950 0.650 2.070 1.850 ;
        RECT  1.640 0.330 1.900 0.500 ;
        RECT  1.705 0.655 1.825 2.140 ;
        RECT  1.465 0.655 1.705 0.775 ;
        RECT  1.225 2.020 1.705 2.140 ;
        RECT  0.945 0.380 1.640 0.500 ;
        RECT  1.225 0.645 1.345 1.630 ;
        RECT  1.070 0.645 1.225 0.815 ;
        RECT  0.810 1.510 1.225 1.630 ;
        RECT  0.985 1.070 1.105 1.390 ;
        RECT  0.255 1.270 0.985 1.390 ;
        RECT  0.825 0.380 0.945 0.740 ;
        RECT  0.230 0.620 0.825 0.740 ;
        RECT  0.230 1.225 0.255 1.555 ;
        RECT  0.085 0.620 0.230 1.555 ;
    END
END CLKMX2X12AD
MACRO CLKMX2X2AD
    CLASS CORE ;
    FOREIGN CLKMX2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.695 0.590 2.730 1.725 ;
        RECT  2.590 0.590 2.695 1.995 ;
        RECT  2.550 0.590 2.590 0.850 ;
        RECT  2.525 1.565 2.590 1.995 ;
        END
        AntennaDiffArea 0.29 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.050 0.230 1.655 ;
        END
        AntennaGateArea 0.1775 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.990 0.780 1.655 ;
        END
        AntennaGateArea 0.1 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.865 2.170 1.375 ;
        END
        AntennaGateArea 0.1 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.360 -0.210 2.800 0.210 ;
        RECT  2.100 -0.210 2.360 0.250 ;
        RECT  0.790 -0.210 2.100 0.210 ;
        RECT  0.530 -0.210 0.790 0.630 ;
        RECT  0.000 -0.210 0.530 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.335 2.310 2.800 2.730 ;
        RECT  2.165 1.565 2.335 2.730 ;
        RECT  0.765 2.310 2.165 2.730 ;
        RECT  0.595 1.815 0.765 2.730 ;
        RECT  0.000 2.310 0.595 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.430 0.990 2.460 1.250 ;
        RECT  2.310 0.550 2.430 1.250 ;
        RECT  2.150 0.550 2.310 0.670 ;
        RECT  2.030 0.400 2.150 0.670 ;
        RECT  1.670 0.400 2.030 0.520 ;
        RECT  1.910 1.540 1.975 1.970 ;
        RECT  1.790 0.640 1.910 1.970 ;
        RECT  1.550 0.400 1.670 1.910 ;
        RECT  1.385 0.400 1.550 0.630 ;
        RECT  1.365 1.740 1.550 1.910 ;
        RECT  1.310 0.750 1.430 1.570 ;
        RECT  1.260 0.750 1.310 0.870 ;
        RECT  1.175 1.450 1.310 1.570 ;
        RECT  1.140 0.510 1.260 0.870 ;
        RECT  1.020 0.990 1.190 1.250 ;
        RECT  1.005 1.450 1.175 1.925 ;
        RECT  0.910 0.510 1.140 0.630 ;
        RECT  0.900 0.750 1.020 1.250 ;
        RECT  0.470 0.750 0.900 0.870 ;
        RECT  0.350 0.750 0.470 1.985 ;
        RECT  0.330 0.750 0.350 0.870 ;
        RECT  0.185 1.815 0.350 1.985 ;
        RECT  0.210 0.500 0.330 0.870 ;
    END
END CLKMX2X2AD
MACRO CLKMX2X3AD
    CLASS CORE ;
    FOREIGN CLKMX2X3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.860 0.525 3.010 1.995 ;
        RECT  2.770 0.525 2.860 0.785 ;
        RECT  2.745 1.735 2.860 1.995 ;
        END
        AntennaDiffArea 0.295 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.030 1.560 1.815 ;
        RECT  0.240 1.695 1.440 1.815 ;
        RECT  0.240 2.050 0.345 2.170 ;
        RECT  0.070 1.695 0.240 2.170 ;
        END
        AntennaGateArea 0.1924 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.800 1.095 ;
        END
        AntennaGateArea 0.126 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.850 2.450 1.300 ;
        END
        AntennaGateArea 0.126 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.555 -0.210 3.360 0.210 ;
        RECT  2.385 -0.210 2.555 0.725 ;
        RECT  0.605 -0.210 2.385 0.210 ;
        RECT  0.435 -0.210 0.605 0.370 ;
        RECT  0.000 -0.210 0.435 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.290 2.310 3.360 2.730 ;
        RECT  3.250 1.780 3.290 2.730 ;
        RECT  3.130 1.570 3.250 2.730 ;
        RECT  2.600 2.310 3.130 2.730 ;
        RECT  2.340 1.900 2.600 2.730 ;
        RECT  0.655 2.310 2.340 2.730 ;
        RECT  0.490 1.945 0.655 2.730 ;
        RECT  0.000 2.310 0.490 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.620 1.005 2.740 1.615 ;
        RECT  2.515 1.495 2.620 1.615 ;
        RECT  2.395 1.495 2.515 1.780 ;
        RECT  1.810 1.660 2.395 1.780 ;
        RECT  2.170 1.400 2.240 1.520 ;
        RECT  2.050 0.630 2.170 1.520 ;
        RECT  1.980 1.400 2.050 1.520 ;
        RECT  1.655 0.330 1.915 0.500 ;
        RECT  1.690 0.665 1.810 2.125 ;
        RECT  1.515 0.665 1.690 0.835 ;
        RECT  1.275 1.955 1.690 2.125 ;
        RECT  0.905 0.380 1.655 0.500 ;
        RECT  1.200 0.635 1.320 1.575 ;
        RECT  1.040 0.635 1.200 0.805 ;
        RECT  0.780 1.455 1.200 1.575 ;
        RECT  0.960 1.020 1.080 1.335 ;
        RECT  0.255 1.215 0.960 1.335 ;
        RECT  0.785 0.380 0.905 0.710 ;
        RECT  0.230 0.590 0.785 0.710 ;
        RECT  0.230 1.215 0.255 1.545 ;
        RECT  0.085 0.590 0.230 1.545 ;
    END
END CLKMX2X3AD
MACRO CLKMX2X4AD
    CLASS CORE ;
    FOREIGN CLKMX2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 0.425 3.010 2.165 ;
        RECT  2.840 0.425 2.870 0.855 ;
        RECT  2.745 1.735 2.870 2.165 ;
        END
        AntennaDiffArea 0.391 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.040 1.560 1.815 ;
        RECT  0.240 1.695 1.440 1.815 ;
        RECT  0.240 2.050 0.345 2.170 ;
        RECT  0.070 1.695 0.240 2.170 ;
        END
        AntennaGateArea 0.1924 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.800 1.095 ;
        END
        AntennaGateArea 0.126 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.850 2.450 1.300 ;
        END
        AntennaGateArea 0.126 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.630 -0.210 3.360 0.210 ;
        RECT  2.460 -0.210 2.630 0.675 ;
        RECT  0.605 -0.210 2.460 0.210 ;
        RECT  0.435 -0.210 0.605 0.370 ;
        RECT  0.000 -0.210 0.435 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.290 2.310 3.360 2.730 ;
        RECT  3.130 1.540 3.290 2.730 ;
        RECT  2.600 2.310 3.130 2.730 ;
        RECT  2.340 1.900 2.600 2.730 ;
        RECT  0.655 2.310 2.340 2.730 ;
        RECT  0.490 1.945 0.655 2.730 ;
        RECT  0.000 2.310 0.490 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.620 1.005 2.740 1.615 ;
        RECT  2.515 1.495 2.620 1.615 ;
        RECT  2.395 1.495 2.515 1.780 ;
        RECT  1.810 1.660 2.395 1.780 ;
        RECT  2.170 1.400 2.240 1.520 ;
        RECT  2.050 0.630 2.170 1.520 ;
        RECT  1.980 1.400 2.050 1.520 ;
        RECT  1.655 0.330 1.915 0.500 ;
        RECT  1.690 0.675 1.810 2.125 ;
        RECT  1.515 0.675 1.690 0.845 ;
        RECT  1.275 1.955 1.690 2.125 ;
        RECT  0.905 0.380 1.655 0.500 ;
        RECT  1.200 0.635 1.320 1.575 ;
        RECT  1.040 0.635 1.200 0.805 ;
        RECT  0.780 1.455 1.200 1.575 ;
        RECT  0.960 1.020 1.080 1.335 ;
        RECT  0.255 1.215 0.960 1.335 ;
        RECT  0.785 0.380 0.905 0.710 ;
        RECT  0.230 0.590 0.785 0.710 ;
        RECT  0.230 1.215 0.255 1.545 ;
        RECT  0.085 0.590 0.230 1.545 ;
    END
END CLKMX2X4AD
MACRO CLKMX2X6AD
    CLASS CORE ;
    FOREIGN CLKMX2X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.600 1.375 3.635 2.065 ;
        RECT  3.430 0.685 3.600 2.065 ;
        RECT  2.915 0.685 3.430 0.855 ;
        RECT  3.010 1.430 3.430 1.550 ;
        RECT  2.860 1.430 3.010 2.165 ;
        RECT  2.745 0.425 2.915 0.855 ;
        RECT  2.745 1.735 2.860 2.165 ;
        END
        AntennaDiffArea 0.584 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.040 1.560 1.815 ;
        RECT  0.240 1.695 1.440 1.815 ;
        RECT  0.240 2.050 0.345 2.170 ;
        RECT  0.070 1.695 0.240 2.170 ;
        END
        AntennaGateArea 0.1924 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.800 1.095 ;
        END
        AntennaGateArea 0.126 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.865 2.450 1.300 ;
        END
        AntennaGateArea 0.126 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.320 -0.210 3.920 0.210 ;
        RECT  3.060 -0.210 3.320 0.550 ;
        RECT  2.555 -0.210 3.060 0.210 ;
        RECT  2.385 -0.210 2.555 0.735 ;
        RECT  0.605 -0.210 2.385 0.210 ;
        RECT  0.435 -0.210 0.605 0.370 ;
        RECT  0.000 -0.210 0.435 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.290 2.310 3.920 2.730 ;
        RECT  3.130 1.670 3.290 2.730 ;
        RECT  2.600 2.310 3.130 2.730 ;
        RECT  2.340 1.900 2.600 2.730 ;
        RECT  0.655 2.310 2.340 2.730 ;
        RECT  0.490 1.945 0.655 2.730 ;
        RECT  0.000 2.310 0.490 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  2.740 1.055 3.165 1.225 ;
        RECT  2.620 1.055 2.740 1.615 ;
        RECT  2.515 1.495 2.620 1.615 ;
        RECT  2.395 1.495 2.515 1.780 ;
        RECT  1.810 1.660 2.395 1.780 ;
        RECT  2.170 1.400 2.240 1.520 ;
        RECT  2.050 0.630 2.170 1.520 ;
        RECT  1.980 1.400 2.050 1.520 ;
        RECT  1.655 0.330 1.915 0.500 ;
        RECT  1.690 0.675 1.810 2.125 ;
        RECT  1.515 0.675 1.690 0.845 ;
        RECT  1.275 1.955 1.690 2.125 ;
        RECT  0.905 0.380 1.655 0.500 ;
        RECT  1.200 0.635 1.320 1.575 ;
        RECT  1.040 0.635 1.200 0.805 ;
        RECT  0.780 1.455 1.200 1.575 ;
        RECT  0.960 1.020 1.080 1.335 ;
        RECT  0.255 1.215 0.960 1.335 ;
        RECT  0.785 0.380 0.905 0.710 ;
        RECT  0.230 0.590 0.785 0.710 ;
        RECT  0.230 1.215 0.255 1.545 ;
        RECT  0.085 0.590 0.230 1.545 ;
    END
END CLKMX2X6AD
MACRO CLKMX2X8AD
    CLASS CORE ;
    FOREIGN CLKMX2X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.635 0.725 3.710 1.470 ;
        RECT  3.465 0.555 3.635 2.065 ;
        RECT  3.290 0.720 3.465 1.470 ;
        RECT  2.915 0.720 3.290 0.890 ;
        RECT  2.985 1.300 3.290 1.470 ;
        RECT  2.865 1.300 2.985 2.165 ;
        RECT  2.745 0.555 2.915 0.890 ;
        RECT  2.745 1.735 2.865 2.165 ;
        END
        AntennaDiffArea 0.699 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.040 1.560 1.815 ;
        RECT  0.240 1.695 1.440 1.815 ;
        RECT  0.240 2.050 0.345 2.170 ;
        RECT  0.070 1.695 0.240 2.170 ;
        END
        AntennaGateArea 0.1924 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.800 1.095 ;
        END
        AntennaGateArea 0.126 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.865 2.450 1.300 ;
        END
        AntennaGateArea 0.126 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.320 -0.210 4.200 0.210 ;
        RECT  3.060 -0.210 3.320 0.600 ;
        RECT  2.555 -0.210 3.060 0.210 ;
        RECT  2.385 -0.210 2.555 0.735 ;
        RECT  0.605 -0.210 2.385 0.210 ;
        RECT  0.435 -0.210 0.605 0.370 ;
        RECT  0.000 -0.210 0.435 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.995 2.310 4.200 2.730 ;
        RECT  3.825 1.585 3.995 2.730 ;
        RECT  3.275 2.310 3.825 2.730 ;
        RECT  3.105 1.595 3.275 2.730 ;
        RECT  2.600 2.310 3.105 2.730 ;
        RECT  2.340 1.900 2.600 2.730 ;
        RECT  0.655 2.310 2.340 2.730 ;
        RECT  0.490 1.945 0.655 2.730 ;
        RECT  0.000 2.310 0.490 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  2.740 1.010 3.165 1.180 ;
        RECT  2.620 1.010 2.740 1.615 ;
        RECT  2.515 1.495 2.620 1.615 ;
        RECT  2.395 1.495 2.515 1.780 ;
        RECT  1.810 1.660 2.395 1.780 ;
        RECT  2.170 1.400 2.240 1.520 ;
        RECT  2.050 0.630 2.170 1.520 ;
        RECT  1.980 1.400 2.050 1.520 ;
        RECT  1.655 0.330 1.915 0.500 ;
        RECT  1.690 0.675 1.810 2.125 ;
        RECT  1.515 0.675 1.690 0.845 ;
        RECT  1.275 1.955 1.690 2.125 ;
        RECT  0.905 0.380 1.655 0.500 ;
        RECT  1.200 0.635 1.320 1.575 ;
        RECT  1.040 0.635 1.200 0.805 ;
        RECT  0.780 1.455 1.200 1.575 ;
        RECT  0.960 1.020 1.080 1.335 ;
        RECT  0.255 1.215 0.960 1.335 ;
        RECT  0.785 0.380 0.905 0.710 ;
        RECT  0.230 0.590 0.785 0.710 ;
        RECT  0.230 1.215 0.255 1.545 ;
        RECT  0.085 0.590 0.230 1.545 ;
    END
END CLKMX2X8AD
MACRO CLKNAND2X12AD
    CLASS CORE ;
    FOREIGN CLKNAND2X12AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.215 0.420 4.660 1.865 ;
        RECT  4.120 0.420 4.215 2.075 ;
        RECT  0.760 0.420 4.120 0.700 ;
        RECT  4.045 1.580 4.120 2.075 ;
        RECT  3.495 1.580 4.045 1.865 ;
        RECT  3.325 1.580 3.495 2.075 ;
        RECT  2.775 1.580 3.325 1.865 ;
        RECT  2.605 1.580 2.775 2.075 ;
        RECT  2.055 1.580 2.605 1.865 ;
        RECT  1.885 1.580 2.055 2.075 ;
        RECT  1.335 1.580 1.885 1.865 ;
        RECT  1.165 1.580 1.335 2.075 ;
        RECT  0.615 1.580 1.165 1.865 ;
        RECT  0.445 1.500 0.615 2.190 ;
        END
        AntennaDiffArea 1.855 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 0.870 3.990 0.990 ;
        RECT  3.160 0.870 3.280 1.170 ;
        RECT  2.810 1.050 3.160 1.170 ;
        RECT  2.690 0.870 2.810 1.170 ;
        RECT  1.860 0.870 2.690 0.990 ;
        RECT  1.340 0.870 1.860 1.170 ;
        RECT  0.490 0.870 1.340 0.990 ;
        RECT  0.320 0.870 0.490 1.375 ;
        END
        AntennaGateArea 0.834 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.540 1.140 3.680 1.260 ;
        RECT  3.420 1.140 3.540 1.410 ;
        RECT  2.470 1.290 3.420 1.410 ;
        RECT  2.210 1.110 2.470 1.410 ;
        RECT  1.140 1.290 2.210 1.410 ;
        RECT  0.910 1.120 1.140 1.410 ;
        RECT  0.620 1.120 0.910 1.375 ;
        END
        AntennaGateArea 0.8349 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.125 -0.210 4.760 0.210 ;
        RECT  2.865 -0.210 3.125 0.300 ;
        RECT  1.740 -0.210 2.865 0.210 ;
        RECT  1.480 -0.210 1.740 0.300 ;
        RECT  0.315 -0.210 1.480 0.210 ;
        RECT  0.145 -0.210 0.315 0.685 ;
        RECT  0.000 -0.210 0.145 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.575 2.310 4.760 2.730 ;
        RECT  4.405 1.985 4.575 2.730 ;
        RECT  3.855 2.310 4.405 2.730 ;
        RECT  3.685 1.985 3.855 2.730 ;
        RECT  3.135 2.310 3.685 2.730 ;
        RECT  2.965 1.985 3.135 2.730 ;
        RECT  2.415 2.310 2.965 2.730 ;
        RECT  2.245 1.985 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 1.985 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.985 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.500 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.760 2.520 ;
	 END
END CLKNAND2X12AD
MACRO CLKNAND2X2AD
    CLASS CORE ;
    FOREIGN CLKNAND2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.585 1.050 1.615 ;
        RECT  0.845 0.585 0.910 0.755 ;
        RECT  0.655 1.495 0.910 1.615 ;
        RECT  0.485 1.495 0.655 1.925 ;
        END
        AntennaDiffArea 0.352 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.240 1.375 ;
        END
        AntennaGateArea 0.141 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 0.875 0.770 1.375 ;
        END
        AntennaGateArea 0.141 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.295 -0.210 1.120 0.210 ;
        RECT  0.125 -0.210 0.295 0.745 ;
        RECT  0.000 -0.210 0.125 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 2.310 1.120 2.730 ;
        RECT  0.845 1.735 1.015 2.730 ;
        RECT  0.295 2.310 0.845 2.730 ;
        RECT  0.125 1.495 0.295 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
	 END
END CLKNAND2X2AD
MACRO CLKNAND2X4AD
    CLASS CORE ;
    FOREIGN CLKNAND2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.715 1.890 1.640 ;
        RECT  1.325 0.715 1.750 0.855 ;
        RECT  1.395 1.500 1.750 1.640 ;
        RECT  1.225 1.500 1.395 2.190 ;
        RECT  1.185 0.555 1.325 0.855 ;
        RECT  0.675 1.500 1.225 1.640 ;
        RECT  0.820 0.555 1.185 0.695 ;
        RECT  0.505 1.500 0.675 2.190 ;
        END
        AntennaDiffArea 0.608 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.040 1.470 1.375 ;
        RECT  0.500 1.255 1.350 1.375 ;
        RECT  0.350 0.865 0.500 1.375 ;
        END
        AntennaGateArea 0.282 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 1.015 1.135 1.135 ;
        RECT  0.630 0.865 0.890 1.135 ;
        END
        AntennaGateArea 0.282 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.645 -0.210 1.960 0.210 ;
        RECT  1.475 -0.210 1.645 0.595 ;
        RECT  0.425 -0.210 1.475 0.210 ;
        RECT  0.255 -0.210 0.425 0.660 ;
        RECT  0.000 -0.210 0.255 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.755 2.310 1.960 2.730 ;
        RECT  1.585 1.845 1.755 2.730 ;
        RECT  1.035 2.310 1.585 2.730 ;
        RECT  0.865 1.845 1.035 2.730 ;
        RECT  0.315 2.310 0.865 2.730 ;
        RECT  0.145 1.585 0.315 2.730 ;
        RECT  0.000 2.310 0.145 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
	 END
END CLKNAND2X4AD
MACRO CLKNAND2X8AD
    CLASS CORE ;
    FOREIGN CLKNAND2X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.030 0.440 3.260 1.820 ;
        RECT  2.460 0.440 3.030 0.670 ;
        RECT  2.775 1.285 3.030 1.820 ;
        RECT  2.730 1.285 2.775 2.075 ;
        RECT  2.605 1.580 2.730 2.075 ;
        RECT  2.055 1.580 2.605 1.820 ;
        RECT  2.200 0.355 2.460 0.735 ;
        RECT  1.020 0.440 2.200 0.670 ;
        RECT  1.885 1.580 2.055 2.075 ;
        RECT  1.335 1.580 1.885 1.820 ;
        RECT  1.165 1.580 1.335 2.075 ;
        RECT  0.615 1.580 1.165 1.820 ;
        RECT  0.760 0.355 1.020 0.735 ;
        RECT  0.445 1.500 0.615 2.190 ;
        END
        AntennaDiffArea 1.216 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.780 0.870 2.900 1.145 ;
        RECT  1.950 0.870 2.780 0.990 ;
        RECT  1.270 0.870 1.950 1.035 ;
        RECT  0.490 0.870 1.270 0.990 ;
        RECT  0.350 0.870 0.490 1.375 ;
        END
        AntennaGateArea 0.564 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.110 2.470 1.230 ;
        RECT  2.190 1.110 2.310 1.410 ;
        RECT  1.375 1.290 2.190 1.410 ;
        RECT  1.030 1.185 1.375 1.410 ;
        RECT  0.770 1.120 1.030 1.410 ;
        END
        AntennaGateArea 0.564 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.090 -0.210 3.360 0.210 ;
        RECT  2.830 -0.210 3.090 0.300 ;
        RECT  1.740 -0.210 2.830 0.210 ;
        RECT  1.480 -0.210 1.740 0.300 ;
        RECT  0.410 -0.210 1.480 0.210 ;
        RECT  0.150 -0.210 0.410 0.735 ;
        RECT  0.000 -0.210 0.150 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.135 2.310 3.360 2.730 ;
        RECT  2.965 1.985 3.135 2.730 ;
        RECT  2.415 2.310 2.965 2.730 ;
        RECT  2.245 1.985 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 1.985 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.945 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.500 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
	 END
END CLKNAND2X8AD
MACRO CLKXOR2X12AD
    CLASS CORE ;
    FOREIGN CLKXOR2X12AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.595 0.655 9.640 1.740 ;
        RECT  9.425 0.475 9.595 1.915 ;
        RECT  8.875 0.655 9.425 1.740 ;
        RECT  8.820 0.655 8.875 2.115 ;
        RECT  8.730 0.470 8.820 2.115 ;
        RECT  8.650 0.470 8.730 0.900 ;
        RECT  8.705 1.360 8.730 2.115 ;
        RECT  8.155 1.360 8.705 1.740 ;
        RECT  7.985 1.360 8.155 2.095 ;
        END
        AntennaDiffArea 0.986 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.110 1.680 1.230 ;
        RECT  1.190 1.110 1.610 1.375 ;
        RECT  0.380 1.110 1.190 1.230 ;
        END
        AntennaGateArea 0.625 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 0.910 2.220 1.330 ;
        END
        AntennaGateArea 0.599 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.955 -0.210 10.080 0.210 ;
        RECT  9.785 -0.210 9.955 0.875 ;
        RECT  9.260 -0.210 9.785 0.210 ;
        RECT  9.000 -0.210 9.260 0.465 ;
        RECT  8.460 -0.210 9.000 0.210 ;
        RECT  8.290 -0.210 8.460 0.875 ;
        RECT  7.680 -0.210 8.290 0.210 ;
        RECT  7.420 -0.210 7.680 0.310 ;
        RECT  6.920 -0.210 7.420 0.210 ;
        RECT  6.660 -0.210 6.920 0.310 ;
        RECT  6.160 -0.210 6.660 0.210 ;
        RECT  5.900 -0.210 6.160 0.310 ;
        RECT  2.195 -0.210 5.900 0.210 ;
        RECT  1.935 -0.210 2.195 0.310 ;
        RECT  1.380 -0.210 1.935 0.210 ;
        RECT  1.120 -0.210 1.380 0.750 ;
        RECT  0.660 -0.210 1.120 0.210 ;
        RECT  0.400 -0.210 0.660 0.750 ;
        RECT  0.000 -0.210 0.400 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.955 2.310 10.080 2.730 ;
        RECT  9.785 1.595 9.955 2.730 ;
        RECT  9.280 2.310 9.785 2.730 ;
        RECT  9.020 1.870 9.280 2.730 ;
        RECT  8.560 2.310 9.020 2.730 ;
        RECT  8.300 1.870 8.560 2.730 ;
        RECT  7.840 2.310 8.300 2.730 ;
        RECT  7.580 2.010 7.840 2.730 ;
        RECT  7.140 2.310 7.580 2.730 ;
        RECT  6.880 1.980 7.140 2.730 ;
        RECT  6.400 2.310 6.880 2.730 ;
        RECT  6.140 2.130 6.400 2.730 ;
        RECT  2.055 2.310 6.140 2.730 ;
        RECT  1.885 1.975 2.055 2.730 ;
        RECT  1.340 2.310 1.885 2.730 ;
        RECT  1.160 1.930 1.340 2.730 ;
        RECT  0.615 2.310 1.160 2.730 ;
        RECT  0.445 1.650 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.080 2.520 ;
        LAYER M1 ;
        RECT  7.750 1.070 8.600 1.190 ;
        RECT  7.630 0.430 7.750 1.860 ;
        RECT  5.520 0.430 7.630 0.550 ;
        RECT  6.760 1.740 7.630 1.860 ;
        RECT  7.380 0.750 7.500 1.620 ;
        RECT  5.780 0.750 7.380 0.870 ;
        RECT  6.470 1.500 7.380 1.620 ;
        RECT  6.020 1.110 7.260 1.230 ;
        RECT  6.640 1.740 6.760 2.010 ;
        RECT  5.630 1.890 6.640 2.010 ;
        RECT  6.350 1.500 6.470 1.720 ;
        RECT  5.230 1.600 6.350 1.720 ;
        RECT  5.900 1.110 6.020 1.470 ;
        RECT  4.240 1.350 5.900 1.470 ;
        RECT  5.660 0.750 5.780 0.980 ;
        RECT  2.605 1.110 5.680 1.230 ;
        RECT  2.945 0.860 5.660 0.980 ;
        RECT  5.400 1.890 5.630 2.140 ;
        RECT  5.400 0.430 5.520 0.740 ;
        RECT  3.090 0.620 5.400 0.740 ;
        RECT  4.940 2.020 5.400 2.140 ;
        RECT  5.110 1.600 5.230 1.860 ;
        RECT  2.940 0.380 5.210 0.500 ;
        RECT  4.510 1.600 5.110 1.720 ;
        RECT  4.680 1.850 4.940 2.140 ;
        RECT  3.835 2.020 4.680 2.140 ;
        RECT  4.390 1.600 4.510 1.860 ;
        RECT  3.980 1.350 4.240 1.900 ;
        RECT  3.520 1.350 3.980 1.470 ;
        RECT  3.665 1.605 3.835 2.140 ;
        RECT  3.115 2.020 3.665 2.140 ;
        RECT  3.260 1.350 3.520 1.900 ;
        RECT  2.730 1.350 3.260 1.470 ;
        RECT  2.945 1.605 3.115 2.140 ;
        RECT  2.775 0.675 2.945 0.980 ;
        RECT  2.820 0.380 2.940 0.555 ;
        RECT  1.670 0.435 2.820 0.555 ;
        RECT  2.610 1.350 2.730 2.175 ;
        RECT  1.695 1.735 2.610 1.855 ;
        RECT  2.485 0.675 2.605 1.230 ;
        RECT  2.355 0.675 2.485 1.615 ;
        RECT  2.200 1.495 2.355 1.615 ;
        RECT  1.525 1.620 1.695 2.050 ;
        RECT  1.550 0.435 1.670 0.990 ;
        RECT  0.950 0.870 1.550 0.990 ;
        RECT  0.975 1.620 1.525 1.740 ;
        RECT  0.805 1.400 0.975 2.135 ;
        RECT  0.830 0.630 0.950 0.990 ;
        RECT  0.230 0.870 0.830 0.990 ;
        RECT  0.255 1.400 0.805 1.520 ;
        RECT  0.230 1.400 0.255 2.130 ;
        RECT  0.110 0.620 0.230 2.130 ;
        RECT  0.085 1.440 0.110 2.130 ;
    END
END CLKXOR2X12AD
MACRO CLKXOR2X1AD
    CLASS CORE ;
    FOREIGN CLKXOR2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 0.610 2.730 2.030 ;
        END
        AntennaDiffArea 0.177 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.380 0.950 1.500 ;
        RECT  0.630 0.740 0.770 1.655 ;
        END
        AntennaGateArea 0.0776 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.030 0.240 1.290 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.1546 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.380 -0.210 2.800 0.210 ;
        RECT  2.120 -0.210 2.380 0.310 ;
        RECT  0.690 -0.210 2.120 0.210 ;
        RECT  0.430 -0.210 0.690 0.260 ;
        RECT  0.000 -0.210 0.430 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.380 2.310 2.800 2.730 ;
        RECT  2.120 1.990 2.380 2.730 ;
        RECT  0.755 2.310 2.120 2.730 ;
        RECT  0.495 2.255 0.755 2.730 ;
        RECT  0.000 2.310 0.495 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.330 0.990 2.450 1.870 ;
        RECT  1.570 1.750 2.330 1.870 ;
        RECT  2.080 0.440 2.200 1.210 ;
        RECT  1.540 0.440 2.080 0.560 ;
        RECT  1.960 0.950 2.080 1.210 ;
        RECT  1.810 1.500 2.000 1.620 ;
        RECT  1.810 0.680 1.960 0.800 ;
        RECT  1.690 0.680 1.810 1.620 ;
        RECT  1.500 1.990 1.760 2.190 ;
        RECT  1.450 0.810 1.570 1.870 ;
        RECT  1.420 0.440 1.540 0.690 ;
        RECT  0.510 1.990 1.500 2.110 ;
        RECT  1.310 0.810 1.450 0.930 ;
        RECT  1.190 0.570 1.420 0.690 ;
        RECT  0.950 0.330 1.300 0.450 ;
        RECT  1.070 0.570 1.190 1.805 ;
        RECT  0.925 0.685 1.070 0.855 ;
        RECT  0.995 1.635 1.070 1.805 ;
        RECT  0.830 0.330 0.950 0.565 ;
        RECT  0.510 0.430 0.830 0.565 ;
        RECT  0.390 0.430 0.510 2.110 ;
        RECT  0.085 0.475 0.390 0.645 ;
        RECT  0.110 1.630 0.390 1.890 ;
    END
END CLKXOR2X1AD
MACRO CLKXOR2X2AD
    CLASS CORE ;
    FOREIGN CLKXOR2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 0.560 2.730 2.045 ;
        END
        AntennaDiffArea 0.29 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.330 0.900 1.450 ;
        RECT  0.630 0.700 0.770 1.450 ;
        END
        AntennaGateArea 0.101 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.240 1.375 ;
        END
        AntennaGateArea 0.1566 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.380 -0.210 2.800 0.210 ;
        RECT  2.120 -0.210 2.380 0.295 ;
        RECT  0.635 -0.210 2.120 0.210 ;
        RECT  0.465 -0.210 0.635 0.255 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.335 2.310 2.800 2.730 ;
        RECT  2.165 2.060 2.335 2.730 ;
        RECT  0.730 2.310 2.165 2.730 ;
        RECT  0.470 2.220 0.730 2.730 ;
        RECT  0.000 2.310 0.470 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.330 0.990 2.450 1.870 ;
        RECT  1.570 1.750 2.330 1.870 ;
        RECT  2.080 0.415 2.200 1.230 ;
        RECT  1.570 0.415 2.080 0.535 ;
        RECT  2.020 0.970 2.080 1.230 ;
        RECT  1.895 0.655 1.955 0.825 ;
        RECT  1.895 1.450 1.955 1.620 ;
        RECT  1.775 0.655 1.895 1.620 ;
        RECT  1.500 1.990 1.760 2.190 ;
        RECT  1.570 0.810 1.620 0.930 ;
        RECT  1.450 0.415 1.570 0.690 ;
        RECT  1.450 0.810 1.570 1.870 ;
        RECT  1.245 1.990 1.500 2.110 ;
        RECT  1.215 0.570 1.450 0.690 ;
        RECT  1.360 0.810 1.450 0.930 ;
        RECT  1.425 1.545 1.450 1.805 ;
        RECT  0.965 0.330 1.310 0.450 ;
        RECT  1.125 1.955 1.245 2.110 ;
        RECT  1.095 0.570 1.215 1.820 ;
        RECT  0.480 1.955 1.125 2.075 ;
        RECT  0.905 0.705 1.095 0.875 ;
        RECT  0.995 1.650 1.095 1.820 ;
        RECT  0.845 0.330 0.965 0.580 ;
        RECT  0.480 0.460 0.845 0.580 ;
        RECT  0.360 0.460 0.480 2.075 ;
        RECT  0.255 0.460 0.360 0.590 ;
        RECT  0.110 1.630 0.360 1.890 ;
        RECT  0.085 0.420 0.255 0.590 ;
    END
END CLKXOR2X2AD
MACRO CLKXOR2X4AD
    CLASS CORE ;
    FOREIGN CLKXOR2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.745 0.415 3.850 1.460 ;
        RECT  3.710 0.415 3.745 2.065 ;
        RECT  3.575 0.415 3.710 0.585 ;
        RECT  3.575 1.305 3.710 2.065 ;
        END
        AntennaDiffArea 0.328 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.090 0.705 1.210 ;
        RECT  0.070 1.090 0.210 1.655 ;
        END
        AntennaGateArea 0.2084 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.865 2.450 1.095 ;
        END
        AntennaGateArea 0.2366 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.090 -0.210 4.200 0.210 ;
        RECT  3.970 -0.210 4.090 0.610 ;
        RECT  3.245 -0.210 3.970 0.210 ;
        RECT  3.245 0.395 3.345 0.565 ;
        RECT  2.985 -0.210 3.245 0.565 ;
        RECT  0.690 -0.210 2.985 0.210 ;
        RECT  2.915 0.395 2.985 0.565 ;
        RECT  0.535 -0.210 0.690 0.665 ;
        RECT  0.000 -0.210 0.535 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.105 2.310 4.200 2.730 ;
        RECT  3.935 1.585 4.105 2.730 ;
        RECT  3.385 2.310 3.935 2.730 ;
        RECT  3.215 1.725 3.385 2.730 ;
        RECT  0.980 2.310 3.215 2.730 ;
        RECT  0.860 2.170 0.980 2.730 ;
        RECT  0.265 2.310 0.860 2.730 ;
        RECT  0.110 1.775 0.265 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  3.330 0.740 3.450 1.105 ;
        RECT  3.310 0.965 3.330 1.105 ;
        RECT  3.190 0.965 3.310 1.590 ;
        RECT  2.260 1.470 3.190 1.590 ;
        RECT  2.690 1.215 3.070 1.335 ;
        RECT  2.690 1.920 2.880 2.190 ;
        RECT  2.570 0.370 2.690 1.335 ;
        RECT  2.620 1.720 2.690 2.190 ;
        RECT  2.430 1.720 2.620 2.140 ;
        RECT  1.970 1.215 2.570 1.335 ;
        RECT  1.245 2.020 2.430 2.140 ;
        RECT  2.180 0.370 2.300 0.745 ;
        RECT  2.140 1.470 2.260 1.875 ;
        RECT  1.730 0.625 2.180 0.745 ;
        RECT  1.565 1.755 2.140 1.875 ;
        RECT  0.945 0.385 1.970 0.505 ;
        RECT  1.850 1.215 1.970 1.635 ;
        RECT  1.710 1.515 1.850 1.635 ;
        RECT  1.610 0.625 1.730 1.395 ;
        RECT  1.565 1.275 1.610 1.395 ;
        RECT  1.445 1.275 1.565 1.875 ;
        RECT  1.285 0.965 1.490 1.085 ;
        RECT  1.395 1.705 1.445 1.875 ;
        RECT  1.115 0.665 1.285 1.545 ;
        RECT  1.125 1.845 1.245 2.140 ;
        RECT  0.945 1.845 1.125 1.965 ;
        RECT  0.825 0.385 0.945 1.965 ;
        RECT  0.330 0.820 0.825 0.940 ;
        RECT  0.450 1.445 0.825 1.965 ;
        RECT  0.210 0.360 0.330 0.940 ;
    END
END CLKXOR2X4AD
MACRO CLKXOR2X8AD
    CLASS CORE ;
    FOREIGN CLKXOR2X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.250 1.355 6.270 1.635 ;
        RECT  6.130 0.640 6.250 2.110 ;
        RECT  5.810 0.640 6.130 1.635 ;
        RECT  5.330 0.640 5.810 0.905 ;
        RECT  5.530 1.355 5.810 1.635 ;
        RECT  5.410 1.355 5.530 2.140 ;
        END
        AntennaDiffArea 0.656 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 0.835 0.870 0.995 ;
        RECT  0.350 0.835 0.490 1.450 ;
        END
        AntennaGateArea 0.4145 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 0.865 1.605 1.025 ;
        RECT  1.190 0.865 1.330 1.375 ;
        END
        AntennaGateArea 0.4155 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.610 -0.210 6.720 0.210 ;
        RECT  6.465 -0.210 6.610 0.940 ;
        RECT  5.940 -0.210 6.465 0.210 ;
        RECT  5.680 -0.210 5.940 0.520 ;
        RECT  5.180 -0.210 5.680 0.210 ;
        RECT  4.920 -0.210 5.180 0.350 ;
        RECT  4.380 -0.210 4.920 0.210 ;
        RECT  4.120 -0.210 4.380 0.350 ;
        RECT  1.340 -0.210 4.120 0.210 ;
        RECT  1.220 -0.210 1.340 0.450 ;
        RECT  0.660 -0.210 1.220 0.210 ;
        RECT  0.400 -0.210 0.660 0.450 ;
        RECT  0.000 -0.210 0.400 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.610 2.310 6.720 2.730 ;
        RECT  6.490 1.420 6.610 2.730 ;
        RECT  5.960 2.310 6.490 2.730 ;
        RECT  5.700 2.010 5.960 2.730 ;
        RECT  5.240 2.310 5.700 2.730 ;
        RECT  4.980 2.130 5.240 2.730 ;
        RECT  4.520 2.310 4.980 2.730 ;
        RECT  4.260 2.130 4.520 2.730 ;
        RECT  1.450 2.310 4.260 2.730 ;
        RECT  1.190 2.290 1.450 2.730 ;
        RECT  0.615 2.310 1.190 2.730 ;
        RECT  0.445 1.845 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.720 2.520 ;
        LAYER M1 ;
        RECT  5.135 1.090 5.670 1.210 ;
        RECT  5.015 0.470 5.135 2.010 ;
        RECT  4.015 0.470 5.015 0.590 ;
        RECT  4.135 1.890 5.015 2.010 ;
        RECT  4.760 0.915 4.880 1.750 ;
        RECT  4.715 0.915 4.760 1.035 ;
        RECT  3.860 1.630 4.760 1.750 ;
        RECT  4.545 0.735 4.715 1.035 ;
        RECT  3.580 1.180 4.640 1.300 ;
        RECT  2.700 0.915 4.545 1.035 ;
        RECT  4.015 1.890 4.135 2.140 ;
        RECT  3.735 0.470 4.015 0.795 ;
        RECT  3.585 1.930 4.015 2.140 ;
        RECT  3.740 1.630 3.860 1.785 ;
        RECT  3.395 1.665 3.740 1.785 ;
        RECT  3.190 0.675 3.735 0.795 ;
        RECT  3.355 0.380 3.615 0.555 ;
        RECT  3.035 2.020 3.585 2.140 ;
        RECT  3.460 1.180 3.580 1.545 ;
        RECT  2.675 1.425 3.460 1.545 ;
        RECT  3.225 1.665 3.395 1.835 ;
        RECT  1.580 0.380 3.355 0.500 ;
        RECT  1.905 1.155 3.280 1.275 ;
        RECT  2.840 0.620 3.190 0.795 ;
        RECT  2.865 1.665 3.035 2.140 ;
        RECT  2.315 2.020 2.865 2.140 ;
        RECT  2.275 0.620 2.840 0.740 ;
        RECT  2.440 0.860 2.700 1.035 ;
        RECT  2.505 1.425 2.675 1.830 ;
        RECT  1.955 1.425 2.505 1.545 ;
        RECT  2.160 1.665 2.315 2.140 ;
        RECT  2.105 0.620 2.275 0.790 ;
        RECT  2.145 1.665 2.160 2.095 ;
        RECT  1.835 1.425 1.955 2.020 ;
        RECT  1.735 0.620 1.905 1.275 ;
        RECT  1.785 1.850 1.835 2.020 ;
        RECT  0.975 1.900 1.785 2.020 ;
        RECT  1.685 1.150 1.735 1.275 ;
        RECT  1.515 1.150 1.685 1.645 ;
        RECT  1.460 0.380 1.580 0.690 ;
        RECT  0.975 0.570 1.460 0.690 ;
        RECT  0.805 0.465 0.975 0.690 ;
        RECT  0.805 1.425 0.975 2.115 ;
        RECT  0.255 0.570 0.805 0.690 ;
        RECT  0.230 1.570 0.805 1.690 ;
        RECT  0.210 0.465 0.255 0.690 ;
        RECT  0.210 1.535 0.230 2.055 ;
        RECT  0.085 0.465 0.210 2.055 ;
    END
END CLKXOR2X8AD
MACRO CMPR42X1AD
    CLASS CORE ;
    FOREIGN CMPR42X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.670 0.650 12.810 1.915 ;
        RECT  12.625 0.650 12.670 0.820 ;
        RECT  12.640 1.395 12.670 1.915 ;
        END
        AntennaDiffArea 0.203 ;
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.625 0.240 0.885 ;
        RECT  0.210 1.455 0.240 1.975 ;
        RECT  0.070 0.625 0.210 1.975 ;
        END
        AntennaDiffArea 0.207 ;
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.955 1.145 11.255 1.375 ;
        END
        AntennaGateArea 0.0994 ;
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.435 0.910 8.555 1.205 ;
        RECT  7.820 0.910 8.435 1.050 ;
        RECT  7.680 0.910 7.820 1.260 ;
        RECT  7.235 1.140 7.680 1.260 ;
        RECT  7.065 1.140 7.235 1.355 ;
        END
        AntennaGateArea 0.2312 ;
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.150 1.420 10.335 1.610 ;
        RECT  10.030 0.660 10.150 1.610 ;
        RECT  9.995 0.660 10.030 0.920 ;
        RECT  9.970 1.420 10.030 1.610 ;
        END
        AntennaDiffArea 0.215 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.945 1.980 8.205 2.185 ;
        RECT  1.655 1.980 7.945 2.100 ;
        RECT  1.145 1.980 1.655 2.170 ;
        END
        AntennaGateArea 0.1864 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.540 1.240 4.380 1.360 ;
        RECT  3.420 1.240 3.540 1.845 ;
        RECT  2.605 1.725 3.420 1.845 ;
        RECT  2.605 1.140 2.745 1.310 ;
        RECT  2.485 1.140 2.605 1.845 ;
        RECT  2.315 1.140 2.485 1.455 ;
        RECT  1.430 1.335 2.315 1.455 ;
        RECT  1.310 1.145 1.430 1.455 ;
        RECT  0.910 1.145 1.310 1.375 ;
        END
        AntennaGateArea 0.3092 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.940 0.870 3.060 1.365 ;
        RECT  2.210 0.870 2.940 0.990 ;
        RECT  1.900 0.870 2.210 1.050 ;
        RECT  1.640 0.870 1.900 1.190 ;
        RECT  0.790 0.870 1.640 0.990 ;
        RECT  0.670 0.870 0.790 1.260 ;
        END
        AntennaGateArea 0.2612 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.520 -0.210 12.880 0.210 ;
        RECT  12.260 -0.210 12.520 0.300 ;
        RECT  11.030 -0.210 12.260 0.210 ;
        RECT  10.510 -0.210 11.030 0.415 ;
        RECT  8.405 -0.210 10.510 0.210 ;
        RECT  8.145 -0.210 8.405 0.300 ;
        RECT  6.680 -0.210 8.145 0.210 ;
        RECT  6.420 -0.210 6.680 0.300 ;
        RECT  4.725 -0.210 6.420 0.210 ;
        RECT  4.465 -0.210 4.725 0.300 ;
        RECT  3.260 -0.210 4.465 0.210 ;
        RECT  3.000 -0.210 3.260 0.510 ;
        RECT  2.085 -0.210 3.000 0.210 ;
        RECT  1.915 -0.210 2.085 0.500 ;
        RECT  0.685 -0.210 1.915 0.210 ;
        RECT  0.425 -0.210 0.685 0.310 ;
        RECT  0.000 -0.210 0.425 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.520 2.310 12.880 2.730 ;
        RECT  12.260 2.220 12.520 2.730 ;
        RECT  10.970 2.310 12.260 2.730 ;
        RECT  10.450 2.220 10.970 2.730 ;
        RECT  8.470 2.310 10.450 2.730 ;
        RECT  8.350 2.145 8.470 2.730 ;
        RECT  6.680 2.310 8.350 2.730 ;
        RECT  6.420 2.220 6.680 2.730 ;
        RECT  4.890 2.310 6.420 2.730 ;
        RECT  4.630 2.220 4.890 2.730 ;
        RECT  3.230 2.310 4.630 2.730 ;
        RECT  2.970 2.220 3.230 2.730 ;
        RECT  2.650 2.310 2.970 2.730 ;
        RECT  2.390 2.220 2.650 2.730 ;
        RECT  2.050 2.310 2.390 2.730 ;
        RECT  1.790 2.220 2.050 2.730 ;
        RECT  0.590 2.310 1.790 2.730 ;
        RECT  0.470 1.750 0.590 2.730 ;
        RECT  0.000 2.310 0.470 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 12.880 2.520 ;
        LAYER M1 ;
        RECT  12.380 1.010 12.530 1.270 ;
        RECT  12.260 0.420 12.380 2.100 ;
        RECT  11.630 0.420 12.260 0.540 ;
        RECT  11.610 1.980 12.260 2.100 ;
        RECT  12.020 0.660 12.140 1.860 ;
        RECT  11.240 0.660 12.020 0.780 ;
        RECT  11.355 1.740 12.020 1.860 ;
        RECT  11.760 1.300 11.880 1.620 ;
        RECT  10.815 1.500 11.760 1.620 ;
        RECT  11.500 1.260 11.640 1.380 ;
        RECT  11.380 0.905 11.500 1.380 ;
        RECT  11.110 0.905 11.380 1.025 ;
        RECT  11.230 1.740 11.355 2.100 ;
        RECT  9.525 1.980 11.230 2.100 ;
        RECT  10.990 0.535 11.110 1.025 ;
        RECT  10.390 0.535 10.990 0.655 ;
        RECT  10.815 0.775 10.860 0.895 ;
        RECT  10.765 0.775 10.815 1.620 ;
        RECT  10.695 0.775 10.765 1.860 ;
        RECT  10.600 0.775 10.695 0.895 ;
        RECT  10.645 1.450 10.695 1.860 ;
        RECT  9.845 1.740 10.645 1.860 ;
        RECT  10.445 1.045 10.565 1.305 ;
        RECT  10.390 1.045 10.445 1.165 ;
        RECT  10.270 0.380 10.390 1.165 ;
        RECT  9.035 0.380 10.270 0.500 ;
        RECT  9.725 0.620 9.850 1.570 ;
        RECT  9.675 1.690 9.845 1.860 ;
        RECT  9.495 0.620 9.725 0.740 ;
        RECT  9.525 1.450 9.725 1.570 ;
        RECT  9.275 1.070 9.605 1.330 ;
        RECT  9.405 1.450 9.525 2.100 ;
        RECT  9.155 0.620 9.275 1.925 ;
        RECT  9.020 1.755 9.155 1.925 ;
        RECT  8.915 0.380 9.035 1.550 ;
        RECT  8.590 0.380 8.915 0.505 ;
        RECT  8.675 0.625 8.795 1.905 ;
        RECT  7.735 1.435 8.675 1.605 ;
        RECT  8.495 0.380 8.590 0.540 ;
        RECT  5.945 0.420 8.495 0.540 ;
        RECT  7.550 1.730 8.075 1.850 ;
        RECT  7.560 0.660 8.000 0.780 ;
        RECT  7.440 0.660 7.560 1.020 ;
        RECT  7.430 1.500 7.550 1.850 ;
        RECT  6.945 0.900 7.440 1.020 ;
        RECT  6.945 1.500 7.430 1.620 ;
        RECT  6.185 0.660 7.320 0.780 ;
        RECT  6.705 1.740 7.310 1.860 ;
        RECT  6.825 0.900 6.945 1.620 ;
        RECT  6.605 1.090 6.825 1.260 ;
        RECT  6.585 1.435 6.705 1.860 ;
        RECT  6.185 1.435 6.585 1.555 ;
        RECT  6.295 1.690 6.465 1.860 ;
        RECT  4.890 1.740 6.295 1.860 ;
        RECT  6.065 0.660 6.185 1.555 ;
        RECT  6.060 1.075 6.065 1.555 ;
        RECT  5.680 1.075 6.060 1.195 ;
        RECT  5.825 0.420 5.945 0.740 ;
        RECT  5.770 1.360 5.890 1.620 ;
        RECT  5.430 0.620 5.825 0.740 ;
        RECT  5.430 1.500 5.770 1.620 ;
        RECT  5.535 0.330 5.705 0.500 ;
        RECT  5.560 0.935 5.680 1.195 ;
        RECT  5.190 0.380 5.535 0.500 ;
        RECT  5.310 0.620 5.430 1.620 ;
        RECT  5.070 0.380 5.190 1.605 ;
        RECT  5.010 0.380 5.070 0.745 ;
        RECT  4.890 0.905 4.950 1.165 ;
        RECT  4.770 0.420 4.890 1.860 ;
        RECT  3.740 0.420 4.770 0.540 ;
        RECT  4.000 1.740 4.770 1.860 ;
        RECT  4.530 0.660 4.650 1.620 ;
        RECT  3.550 0.660 4.530 0.780 ;
        RECT  3.780 1.500 4.530 1.620 ;
        RECT  3.300 0.940 4.140 1.060 ;
        RECT  3.660 1.500 3.780 1.760 ;
        RECT  3.430 0.445 3.550 0.780 ;
        RECT  3.180 0.630 3.300 1.605 ;
        RECT  2.815 0.630 3.180 0.750 ;
        RECT  2.770 1.485 3.180 1.605 ;
        RECT  2.645 0.570 2.815 0.750 ;
        RECT  1.475 0.620 2.510 0.740 ;
        RECT  1.465 1.575 2.295 1.745 ;
        RECT  0.490 0.620 1.340 0.740 ;
        RECT  0.825 1.595 1.320 1.715 ;
        RECT  0.705 1.460 0.825 1.715 ;
        RECT  0.490 1.460 0.705 1.580 ;
        RECT  0.370 0.620 0.490 1.580 ;
    END
END CMPR42X1AD
MACRO CMPR42X2AD
    CLASS CORE ;
    FOREIGN CMPR42X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.670 0.330 12.810 2.190 ;
        RECT  12.640 0.330 12.670 0.850 ;
        RECT  12.640 1.410 12.670 2.190 ;
        END
        AntennaDiffArea 0.363 ;
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.625 0.240 0.885 ;
        RECT  0.210 1.410 0.240 2.190 ;
        RECT  0.070 0.625 0.210 2.190 ;
        END
        AntennaDiffArea 0.373 ;
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.955 1.140 11.250 1.375 ;
        END
        AntennaGateArea 0.135 ;
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.435 0.890 8.555 1.205 ;
        RECT  7.810 0.890 8.435 1.050 ;
        RECT  7.690 0.890 7.810 1.240 ;
        RECT  7.235 1.120 7.690 1.240 ;
        RECT  7.065 1.120 7.235 1.365 ;
        END
        AntennaGateArea 0.2925 ;
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.150 1.375 10.335 1.635 ;
        RECT  10.030 0.630 10.150 1.635 ;
        RECT  9.995 0.630 10.030 0.890 ;
        RECT  9.970 1.375 10.030 1.635 ;
        END
        AntennaDiffArea 0.304 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.950 1.980 7.985 2.100 ;
        RECT  7.690 1.980 7.950 2.190 ;
        RECT  1.530 1.980 7.690 2.100 ;
        RECT  1.145 1.980 1.530 2.190 ;
        END
        AntennaGateArea 0.2814 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 1.240 4.390 1.360 ;
        RECT  3.540 1.140 3.760 1.360 ;
        RECT  3.500 1.140 3.540 1.845 ;
        RECT  3.420 1.240 3.500 1.845 ;
        RECT  2.605 1.725 3.420 1.845 ;
        RECT  2.605 1.140 2.745 1.310 ;
        RECT  2.485 1.140 2.605 1.845 ;
        RECT  2.315 1.140 2.485 1.455 ;
        RECT  1.370 1.335 2.315 1.455 ;
        RECT  1.250 1.090 1.370 1.455 ;
        RECT  0.910 1.090 1.250 1.375 ;
        END
        AntennaGateArea 0.4646 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.940 0.850 3.060 1.270 ;
        RECT  2.210 0.850 2.940 0.990 ;
        RECT  1.960 0.850 2.210 1.050 ;
        RECT  1.700 0.850 1.960 1.145 ;
        RECT  0.790 0.850 1.700 0.970 ;
        RECT  0.670 0.850 0.790 1.260 ;
        END
        AntennaGateArea 0.4208 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.435 -0.210 12.880 0.210 ;
        RECT  12.265 -0.210 12.435 0.580 ;
        RECT  10.955 -0.210 12.265 0.210 ;
        RECT  10.525 -0.210 10.955 0.405 ;
        RECT  8.405 -0.210 10.525 0.210 ;
        RECT  8.145 -0.210 8.405 0.270 ;
        RECT  6.580 -0.210 8.145 0.210 ;
        RECT  6.320 -0.210 6.580 0.270 ;
        RECT  4.725 -0.210 6.320 0.210 ;
        RECT  4.465 -0.210 4.725 0.300 ;
        RECT  3.215 -0.210 4.465 0.210 ;
        RECT  3.045 -0.210 3.215 0.490 ;
        RECT  2.130 -0.210 3.045 0.210 ;
        RECT  1.870 -0.210 2.130 0.395 ;
        RECT  0.670 -0.210 1.870 0.210 ;
        RECT  0.410 -0.210 0.670 0.395 ;
        RECT  0.000 -0.210 0.410 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.460 2.310 12.880 2.730 ;
        RECT  12.200 2.290 12.460 2.730 ;
        RECT  10.955 2.310 12.200 2.730 ;
        RECT  10.435 2.235 10.955 2.730 ;
        RECT  8.455 2.310 10.435 2.730 ;
        RECT  8.285 1.740 8.455 2.730 ;
        RECT  6.680 2.310 8.285 2.730 ;
        RECT  6.420 2.220 6.680 2.730 ;
        RECT  4.845 2.310 6.420 2.730 ;
        RECT  4.675 2.220 4.845 2.730 ;
        RECT  3.230 2.310 4.675 2.730 ;
        RECT  2.970 2.220 3.230 2.730 ;
        RECT  2.730 2.310 2.970 2.730 ;
        RECT  2.470 2.220 2.730 2.730 ;
        RECT  1.970 2.310 2.470 2.730 ;
        RECT  1.710 2.220 1.970 2.730 ;
        RECT  0.590 2.310 1.710 2.730 ;
        RECT  0.470 1.750 0.590 2.730 ;
        RECT  0.000 2.310 0.470 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 12.880 2.520 ;
        LAYER M1 ;
        RECT  12.400 0.700 12.520 2.140 ;
        RECT  11.980 0.700 12.400 0.820 ;
        RECT  11.570 2.020 12.400 2.140 ;
        RECT  12.100 0.940 12.220 1.900 ;
        RECT  11.740 0.940 12.100 1.060 ;
        RECT  11.330 1.780 12.100 1.900 ;
        RECT  11.860 0.420 11.980 0.820 ;
        RECT  11.790 1.200 11.910 1.660 ;
        RECT  11.610 0.420 11.860 0.540 ;
        RECT  10.815 1.540 11.790 1.660 ;
        RECT  11.620 0.660 11.740 1.060 ;
        RECT  11.500 1.300 11.650 1.420 ;
        RECT  11.230 0.660 11.620 0.780 ;
        RECT  11.380 0.900 11.500 1.420 ;
        RECT  11.100 0.900 11.380 1.020 ;
        RECT  11.210 1.780 11.330 2.115 ;
        RECT  9.525 1.995 11.210 2.115 ;
        RECT  10.980 0.535 11.100 1.020 ;
        RECT  10.390 0.535 10.980 0.655 ;
        RECT  10.735 0.775 10.815 1.660 ;
        RECT  10.695 0.775 10.735 1.875 ;
        RECT  10.645 0.775 10.695 0.945 ;
        RECT  10.615 1.450 10.695 1.875 ;
        RECT  9.845 1.755 10.615 1.875 ;
        RECT  10.445 1.045 10.565 1.305 ;
        RECT  10.390 1.045 10.445 1.165 ;
        RECT  10.270 0.390 10.390 1.165 ;
        RECT  9.950 0.390 10.270 0.510 ;
        RECT  9.780 0.330 9.950 0.510 ;
        RECT  9.725 0.630 9.845 1.570 ;
        RECT  9.675 1.690 9.845 1.875 ;
        RECT  9.035 0.390 9.780 0.510 ;
        RECT  9.535 0.630 9.725 0.750 ;
        RECT  9.525 1.450 9.725 1.570 ;
        RECT  9.485 1.040 9.605 1.330 ;
        RECT  9.405 1.450 9.525 2.115 ;
        RECT  9.275 1.070 9.485 1.330 ;
        RECT  9.155 0.630 9.275 2.145 ;
        RECT  9.020 1.715 9.155 2.145 ;
        RECT  8.915 0.390 9.035 1.460 ;
        RECT  5.945 0.390 8.915 0.510 ;
        RECT  8.675 0.630 8.795 2.190 ;
        RECT  7.880 1.500 8.675 1.620 ;
        RECT  7.550 1.740 8.075 1.860 ;
        RECT  7.560 0.650 8.000 0.770 ;
        RECT  7.760 1.360 7.880 1.620 ;
        RECT  7.440 0.650 7.560 1.000 ;
        RECT  7.430 1.500 7.550 1.860 ;
        RECT  6.945 0.880 7.440 1.000 ;
        RECT  6.945 1.500 7.430 1.620 ;
        RECT  6.185 0.640 7.320 0.760 ;
        RECT  6.705 1.740 7.310 1.860 ;
        RECT  6.825 0.880 6.945 1.620 ;
        RECT  6.555 1.065 6.825 1.235 ;
        RECT  6.585 1.435 6.705 1.860 ;
        RECT  6.185 1.435 6.585 1.555 ;
        RECT  6.295 1.690 6.465 1.860 ;
        RECT  4.890 1.740 6.295 1.860 ;
        RECT  6.065 0.640 6.185 1.555 ;
        RECT  6.060 1.075 6.065 1.555 ;
        RECT  5.680 1.075 6.060 1.195 ;
        RECT  5.825 0.390 5.945 0.740 ;
        RECT  5.770 1.360 5.890 1.620 ;
        RECT  5.440 0.620 5.825 0.740 ;
        RECT  5.440 1.360 5.770 1.480 ;
        RECT  5.535 0.330 5.705 0.500 ;
        RECT  5.560 0.935 5.680 1.195 ;
        RECT  5.200 0.380 5.535 0.500 ;
        RECT  5.320 0.620 5.440 1.480 ;
        RECT  5.080 0.380 5.200 1.605 ;
        RECT  5.010 0.380 5.080 0.745 ;
        RECT  4.890 0.995 4.950 1.255 ;
        RECT  4.770 0.420 4.890 1.860 ;
        RECT  3.740 0.420 4.770 0.540 ;
        RECT  4.000 1.740 4.770 1.860 ;
        RECT  4.530 0.660 4.650 1.620 ;
        RECT  3.550 0.660 4.530 0.780 ;
        RECT  3.780 1.500 4.530 1.620 ;
        RECT  3.890 0.900 4.150 1.060 ;
        RECT  3.300 0.900 3.890 1.020 ;
        RECT  3.660 1.500 3.780 1.760 ;
        RECT  3.430 0.445 3.550 0.780 ;
        RECT  3.180 0.610 3.300 1.605 ;
        RECT  2.880 0.610 3.180 0.730 ;
        RECT  2.770 1.485 3.180 1.605 ;
        RECT  2.760 0.345 2.880 0.730 ;
        RECT  2.620 0.345 2.760 0.465 ;
        RECT  2.320 0.375 2.440 0.635 ;
        RECT  1.680 0.515 2.320 0.635 ;
        RECT  1.505 1.575 2.305 1.745 ;
        RECT  1.510 0.465 1.680 0.635 ;
        RECT  0.825 1.595 1.310 1.715 ;
        RECT  1.105 0.465 1.275 0.635 ;
        RECT  0.490 0.515 1.105 0.635 ;
        RECT  0.705 1.460 0.825 1.715 ;
        RECT  0.490 1.460 0.705 1.580 ;
        RECT  0.370 0.515 0.490 1.580 ;
    END
END CMPR42X2AD
MACRO CMPR42X4AD
    CLASS CORE ;
    FOREIGN CMPR42X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  18.010 0.615 18.130 1.770 ;
        RECT  17.990 0.355 18.010 2.030 ;
        RECT  17.890 0.355 17.990 0.875 ;
        RECT  17.890 1.510 17.990 2.030 ;
        END
        AntennaDiffArea 0.417 ;
    END S
    PIN ICO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 0.365 0.615 0.795 ;
        RECT  0.490 1.410 0.590 2.190 ;
        RECT  0.470 0.365 0.490 2.190 ;
        RECT  0.350 0.365 0.470 1.780 ;
        END
        AntennaDiffArea 0.422 ;
    END ICO
    PIN ICI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.910 1.140 15.330 1.375 ;
        END
        AntennaGateArea 0.1589 ;
    END ICI
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.775 0.910 10.895 1.240 ;
        RECT  10.390 0.910 10.775 1.100 ;
        RECT  10.105 0.980 10.390 1.100 ;
        RECT  9.985 0.980 10.105 1.280 ;
        RECT  9.675 1.160 9.985 1.280 ;
        RECT  9.415 1.160 9.675 1.310 ;
        END
        AntennaGateArea 0.304 ;
    END D
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.070 0.680 14.210 1.600 ;
        RECT  13.780 0.680 14.070 0.850 ;
        RECT  13.930 1.340 14.070 1.600 ;
        END
        AntennaDiffArea 0.41 ;
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.615 1.980 11.055 2.100 ;
        RECT  10.105 1.980 10.615 2.170 ;
        RECT  8.985 1.980 10.105 2.100 ;
        RECT  8.865 1.980 8.985 2.140 ;
        RECT  8.565 2.020 8.865 2.140 ;
        RECT  8.445 1.980 8.565 2.140 ;
        RECT  3.120 1.980 8.445 2.100 ;
        RECT  3.000 1.980 3.120 2.190 ;
        RECT  2.645 2.070 3.000 2.190 ;
        END
        AntennaGateArea 0.38 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.465 1.220 6.725 1.380 ;
        RECT  6.005 1.260 6.465 1.380 ;
        RECT  5.785 1.140 6.005 1.380 ;
        RECT  5.665 1.140 5.785 1.845 ;
        RECT  4.840 1.725 5.665 1.845 ;
        RECT  4.720 1.140 4.840 1.845 ;
        RECT  4.005 1.140 4.720 1.260 ;
        RECT  3.885 1.140 4.005 1.410 ;
        RECT  1.670 1.290 3.885 1.410 ;
        RECT  1.425 1.175 1.670 1.610 ;
        RECT  1.290 1.175 1.425 1.435 ;
        END
        AntennaGateArea 0.7182 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.065 0.900 5.305 1.365 ;
        RECT  3.765 0.900 5.065 1.020 ;
        RECT  3.645 0.900 3.765 1.170 ;
        RECT  1.920 1.050 3.645 1.170 ;
        RECT  1.800 0.935 1.920 1.170 ;
        RECT  1.100 0.935 1.800 1.055 ;
        RECT  0.980 0.935 1.100 1.260 ;
        END
        AntennaGateArea 0.6818 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.400 -0.210 18.480 0.210 ;
        RECT  18.250 -0.210 18.400 0.885 ;
        RECT  17.700 -0.210 18.250 0.210 ;
        RECT  17.440 -0.210 17.700 0.300 ;
        RECT  16.440 -0.210 17.440 0.210 ;
        RECT  16.180 -0.210 16.440 0.300 ;
        RECT  15.025 -0.210 16.180 0.210 ;
        RECT  14.855 -0.210 15.025 0.300 ;
        RECT  14.375 -0.210 14.855 0.210 ;
        RECT  14.115 -0.210 14.375 0.300 ;
        RECT  13.615 -0.210 14.115 0.210 ;
        RECT  13.355 -0.210 13.615 0.300 ;
        RECT  10.795 -0.210 13.355 0.210 ;
        RECT  10.535 -0.210 10.795 0.260 ;
        RECT  8.925 -0.210 10.535 0.210 ;
        RECT  8.665 -0.210 8.925 0.260 ;
        RECT  6.995 -0.210 8.665 0.210 ;
        RECT  6.735 -0.210 6.995 0.300 ;
        RECT  5.450 -0.210 6.735 0.210 ;
        RECT  5.280 -0.210 5.450 0.540 ;
        RECT  4.345 -0.210 5.280 0.210 ;
        RECT  4.085 -0.210 4.345 0.540 ;
        RECT  3.625 -0.210 4.085 0.210 ;
        RECT  3.365 -0.210 3.625 0.540 ;
        RECT  2.220 -0.210 3.365 0.210 ;
        RECT  2.050 -0.210 2.220 0.340 ;
        RECT  0.975 -0.210 2.050 0.210 ;
        RECT  0.805 -0.210 0.975 0.575 ;
        RECT  0.230 -0.210 0.805 0.210 ;
        RECT  0.085 -0.210 0.230 0.840 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.395 2.310 18.480 2.730 ;
        RECT  18.250 1.435 18.395 2.730 ;
        RECT  17.700 2.310 18.250 2.730 ;
        RECT  17.440 2.220 17.700 2.730 ;
        RECT  16.440 2.310 17.440 2.730 ;
        RECT  16.180 2.220 16.440 2.730 ;
        RECT  14.785 2.310 16.180 2.730 ;
        RECT  14.615 2.265 14.785 2.730 ;
        RECT  13.760 2.310 14.615 2.730 ;
        RECT  13.500 2.220 13.760 2.730 ;
        RECT  11.295 2.310 13.500 2.730 ;
        RECT  11.175 1.640 11.295 2.730 ;
        RECT  10.705 1.640 11.175 1.810 ;
        RECT  8.995 2.310 11.175 2.730 ;
        RECT  8.735 2.260 8.995 2.730 ;
        RECT  7.225 2.310 8.735 2.730 ;
        RECT  6.965 2.220 7.225 2.730 ;
        RECT  5.245 2.310 6.965 2.730 ;
        RECT  4.725 2.220 5.245 2.730 ;
        RECT  3.605 2.310 4.725 2.730 ;
        RECT  3.435 2.265 3.605 2.730 ;
        RECT  2.220 2.310 3.435 2.730 ;
        RECT  2.050 2.105 2.220 2.730 ;
        RECT  0.975 2.310 2.050 2.730 ;
        RECT  0.805 1.795 0.975 2.730 ;
        RECT  0.230 2.310 0.805 2.730 ;
        RECT  0.090 1.440 0.230 2.730 ;
        RECT  0.000 2.310 0.090 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 18.480 2.520 ;
        LAYER M1 ;
        RECT  17.770 0.995 17.860 1.255 ;
        RECT  17.650 0.420 17.770 2.100 ;
        RECT  15.550 0.420 17.650 0.540 ;
        RECT  15.550 1.980 17.650 2.100 ;
        RECT  17.340 0.660 17.460 1.860 ;
        RECT  15.405 0.660 17.340 0.780 ;
        RECT  16.410 1.140 17.340 1.260 ;
        RECT  15.405 1.740 17.340 1.860 ;
        RECT  16.820 1.380 17.080 1.620 ;
        RECT  15.905 0.900 17.070 1.020 ;
        RECT  16.280 1.500 16.820 1.620 ;
        RECT  16.160 1.180 16.280 1.620 ;
        RECT  14.775 1.500 16.160 1.620 ;
        RECT  15.475 0.900 15.905 1.380 ;
        RECT  15.015 0.900 15.475 1.020 ;
        RECT  15.235 0.505 15.405 0.780 ;
        RECT  15.235 1.740 15.405 2.080 ;
        RECT  13.520 1.960 15.235 2.080 ;
        RECT  14.895 0.420 15.015 1.020 ;
        RECT  14.510 0.420 14.895 0.540 ;
        RECT  14.655 0.660 14.775 1.840 ;
        RECT  14.630 0.660 14.655 0.920 ;
        RECT  14.630 1.395 14.655 1.840 ;
        RECT  13.760 1.720 14.630 1.840 ;
        RECT  14.510 1.020 14.535 1.280 ;
        RECT  14.390 0.420 14.510 1.280 ;
        RECT  13.120 0.420 14.390 0.540 ;
        RECT  13.640 1.430 13.760 1.840 ;
        RECT  13.330 1.430 13.640 1.550 ;
        RECT  13.400 1.675 13.520 2.080 ;
        RECT  13.365 0.660 13.485 1.260 ;
        RECT  13.210 1.675 13.400 1.795 ;
        RECT  12.855 0.660 13.365 0.780 ;
        RECT  13.210 1.140 13.365 1.260 ;
        RECT  13.160 1.915 13.280 2.175 ;
        RECT  12.970 0.900 13.245 1.020 ;
        RECT  13.090 1.140 13.210 1.795 ;
        RECT  12.585 2.020 13.160 2.140 ;
        RECT  13.000 0.380 13.120 0.540 ;
        RECT  12.945 1.675 13.090 1.795 ;
        RECT  12.275 0.380 13.000 0.500 ;
        RECT  12.850 0.900 12.970 1.270 ;
        RECT  12.775 1.675 12.945 1.845 ;
        RECT  12.595 0.620 12.855 0.780 ;
        RECT  12.585 1.050 12.850 1.270 ;
        RECT  12.450 1.050 12.585 2.140 ;
        RECT  12.355 0.620 12.475 0.740 ;
        RECT  12.355 1.050 12.450 1.170 ;
        RECT  11.775 1.970 12.450 2.140 ;
        RECT  12.235 0.620 12.355 1.170 ;
        RECT  12.050 1.605 12.305 1.775 ;
        RECT  12.015 0.330 12.275 0.500 ;
        RECT  11.635 0.620 12.235 0.740 ;
        RECT  12.050 0.860 12.115 0.980 ;
        RECT  11.920 0.860 12.050 1.775 ;
        RECT  11.395 0.380 12.015 0.500 ;
        RECT  11.855 0.860 11.920 0.980 ;
        RECT  11.585 1.650 11.920 1.775 ;
        RECT  11.680 1.160 11.800 1.520 ;
        RECT  11.395 1.160 11.680 1.280 ;
        RECT  11.515 0.620 11.635 0.880 ;
        RECT  11.535 1.650 11.585 2.100 ;
        RECT  11.415 1.400 11.535 2.100 ;
        RECT  11.155 1.400 11.415 1.520 ;
        RECT  11.275 0.380 11.395 1.280 ;
        RECT  8.280 0.380 11.275 0.500 ;
        RECT  11.035 0.625 11.155 1.520 ;
        RECT  10.055 1.400 11.035 1.520 ;
        RECT  9.915 1.690 10.400 1.860 ;
        RECT  9.860 0.660 10.365 0.780 ;
        RECT  9.795 1.500 9.915 1.860 ;
        RECT  9.740 0.660 9.860 1.030 ;
        RECT  9.295 1.500 9.795 1.620 ;
        RECT  9.295 0.910 9.740 1.030 ;
        RECT  9.055 1.740 9.675 1.860 ;
        RECT  8.565 0.630 9.620 0.750 ;
        RECT  9.175 0.910 9.295 1.620 ;
        RECT  8.850 1.025 9.175 1.195 ;
        RECT  8.935 1.400 9.055 1.860 ;
        RECT  8.565 1.400 8.935 1.520 ;
        RECT  8.655 1.640 8.775 1.900 ;
        RECT  7.225 1.740 8.655 1.860 ;
        RECT  8.445 0.630 8.565 1.520 ;
        RECT  8.395 1.030 8.445 1.520 ;
        RECT  8.075 1.030 8.395 1.150 ;
        RECT  8.160 0.380 8.280 0.810 ;
        RECT  8.080 1.450 8.250 1.620 ;
        RECT  7.775 0.690 8.160 0.810 ;
        RECT  7.775 1.450 8.080 1.570 ;
        RECT  7.955 1.030 8.075 1.290 ;
        RECT  7.870 0.355 8.040 0.525 ;
        RECT  7.535 0.405 7.870 0.525 ;
        RECT  7.655 0.690 7.775 1.570 ;
        RECT  7.415 0.405 7.535 1.620 ;
        RECT  7.345 0.405 7.415 0.745 ;
        RECT  7.225 1.000 7.285 1.260 ;
        RECT  7.105 0.420 7.225 1.860 ;
        RECT  5.985 0.420 7.105 0.540 ;
        RECT  6.285 1.740 7.105 1.860 ;
        RECT  6.865 0.660 6.985 1.620 ;
        RECT  5.810 0.660 6.865 0.780 ;
        RECT  6.025 1.500 6.865 1.620 ;
        RECT  6.125 0.900 6.385 1.130 ;
        RECT  5.545 0.900 6.125 1.020 ;
        RECT  5.905 1.500 6.025 1.760 ;
        RECT  5.690 0.395 5.810 0.780 ;
        RECT  5.640 0.395 5.690 0.565 ;
        RECT  5.425 0.660 5.545 1.605 ;
        RECT  5.045 0.660 5.425 0.780 ;
        RECT  5.025 1.485 5.425 1.605 ;
        RECT  4.925 0.505 5.045 0.780 ;
        RECT  4.515 0.505 4.635 0.780 ;
        RECT  3.220 1.625 4.600 1.795 ;
        RECT  3.220 0.660 4.515 0.780 ;
        RECT  3.050 0.510 3.220 0.780 ;
        RECT  3.050 1.530 3.220 1.795 ;
        RECT  2.285 0.510 3.050 0.630 ;
        RECT  2.285 1.530 3.050 1.650 ;
        RECT  2.165 0.750 2.905 0.870 ;
        RECT  1.585 1.770 2.905 1.890 ;
        RECT  2.040 0.695 2.165 0.870 ;
        RECT  1.590 0.695 2.040 0.815 ;
        RECT  1.420 0.560 1.590 0.815 ;
        RECT  1.415 1.730 1.585 2.160 ;
        RECT  0.855 0.695 1.420 0.815 ;
        RECT  1.255 1.730 1.415 1.890 ;
        RECT  1.135 1.555 1.255 1.890 ;
        RECT  0.855 1.555 1.135 1.675 ;
        RECT  0.735 0.695 0.855 1.675 ;
        RECT  0.620 1.020 0.735 1.280 ;
    END
END CMPR42X4AD
MACRO DFFHQX1AD
    CLASS CORE ;
    FOREIGN DFFHQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.300 0.865 6.370 1.375 ;
        RECT  6.250 0.420 6.300 1.950 ;
        RECT  6.160 0.420 6.250 1.995 ;
        RECT  6.030 0.420 6.160 0.540 ;
        RECT  6.130 1.735 6.160 1.995 ;
        END
        AntennaDiffArea 0.219 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.000 1.890 1.260 ;
        RECT  1.610 1.100 1.770 1.260 ;
        RECT  1.470 1.100 1.610 1.375 ;
        END
        AntennaGateArea 0.077 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.170 1.715 0.535 1.890 ;
        END
        AntennaGateArea 0.114 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.635 -0.210 6.720 0.210 ;
        RECT  6.490 -0.210 6.635 0.915 ;
        RECT  5.695 -0.210 6.490 0.210 ;
        RECT  5.435 -0.210 5.695 0.370 ;
        RECT  3.850 -0.210 5.435 0.210 ;
        RECT  3.590 -0.210 3.850 0.300 ;
        RECT  2.460 -0.210 3.590 0.210 ;
        RECT  2.200 -0.210 2.460 0.300 ;
        RECT  1.765 -0.210 2.200 0.210 ;
        RECT  1.505 -0.210 1.765 0.300 ;
        RECT  0.600 -0.210 1.505 0.210 ;
        RECT  0.600 0.750 0.670 0.870 ;
        RECT  0.480 -0.210 0.600 0.870 ;
        RECT  0.000 -0.210 0.480 0.210 ;
        RECT  0.410 0.750 0.480 0.870 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.635 2.310 6.720 2.730 ;
        RECT  6.465 1.460 6.635 2.730 ;
        RECT  5.660 2.310 6.465 2.730 ;
        RECT  5.400 2.180 5.660 2.730 ;
        RECT  4.125 2.310 5.400 2.730 ;
        RECT  3.605 2.220 4.125 2.730 ;
        RECT  2.490 2.310 3.605 2.730 ;
        RECT  2.230 2.220 2.490 2.730 ;
        RECT  1.890 2.310 2.230 2.730 ;
        RECT  1.630 2.220 1.890 2.730 ;
        RECT  0.600 2.310 1.630 2.730 ;
        RECT  0.340 2.010 0.600 2.730 ;
        RECT  0.000 2.310 0.340 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.720 2.520 ;
        LAYER M1 ;
        RECT  5.850 0.690 5.970 1.590 ;
        RECT  5.720 1.905 5.920 2.025 ;
        RECT  5.480 1.120 5.850 1.240 ;
        RECT  5.600 1.700 5.720 2.025 ;
        RECT  4.870 1.700 5.600 1.820 ;
        RECT  5.360 0.980 5.480 1.240 ;
        RECT  5.020 0.380 5.140 1.370 ;
        RECT  4.860 1.960 5.120 2.190 ;
        RECT  5.000 0.380 5.020 0.500 ;
        RECT  4.740 0.330 5.000 0.500 ;
        RECT  4.870 0.630 4.900 0.750 ;
        RECT  4.750 0.630 4.870 1.820 ;
        RECT  1.625 1.960 4.860 2.080 ;
        RECT  4.640 0.630 4.750 0.750 ;
        RECT  4.060 0.380 4.740 0.500 ;
        RECT  4.465 1.400 4.515 1.830 ;
        RECT  4.345 0.630 4.465 1.830 ;
        RECT  4.170 0.630 4.345 0.750 ;
        RECT  2.510 1.710 4.345 1.830 ;
        RECT  4.090 0.880 4.210 1.590 ;
        RECT  3.430 1.470 4.090 1.590 ;
        RECT  3.940 0.380 4.060 0.540 ;
        RECT  3.670 0.420 3.940 0.540 ;
        RECT  3.550 0.420 3.670 1.340 ;
        RECT  2.960 0.420 3.550 0.540 ;
        RECT  3.310 0.710 3.430 1.590 ;
        RECT  2.870 0.710 3.310 0.830 ;
        RECT  2.920 1.440 3.310 1.590 ;
        RECT  3.070 0.990 3.190 1.250 ;
        RECT  2.750 0.990 3.070 1.110 ;
        RECT  2.700 0.370 2.960 0.540 ;
        RECT  2.630 0.680 2.750 1.110 ;
        RECT  0.960 0.420 2.700 0.540 ;
        RECT  2.130 0.680 2.630 0.800 ;
        RECT  2.390 0.970 2.510 1.830 ;
        RECT  2.010 0.680 2.130 1.590 ;
        RECT  1.850 0.680 2.010 0.850 ;
        RECT  1.505 1.710 1.625 2.080 ;
        RECT  1.270 1.710 1.505 1.830 ;
        RECT  1.120 1.950 1.380 2.170 ;
        RECT  1.270 0.675 1.335 0.845 ;
        RECT  1.150 0.675 1.270 1.830 ;
        RECT  1.060 1.415 1.150 1.675 ;
        RECT  0.990 1.950 1.120 2.070 ;
        RECT  0.930 1.845 0.990 2.070 ;
        RECT  0.930 0.420 0.960 0.920 ;
        RECT  0.810 0.420 0.930 2.070 ;
        RECT  0.775 1.845 0.810 2.070 ;
        RECT  0.730 1.845 0.775 1.965 ;
        RECT  0.570 0.990 0.690 1.250 ;
        RECT  0.265 1.060 0.570 1.180 ;
        RECT  0.240 0.815 0.265 1.595 ;
        RECT  0.145 0.680 0.240 1.595 ;
        RECT  0.120 0.680 0.145 0.940 ;
        RECT  0.120 1.335 0.145 1.595 ;
    END
END DFFHQX1AD
MACRO DFFHQX2AD
    CLASS CORE ;
    FOREIGN DFFHQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.890 0.685 6.930 1.580 ;
        RECT  6.790 0.355 6.890 2.170 ;
        RECT  6.730 0.355 6.790 0.875 ;
        RECT  6.730 1.390 6.790 2.170 ;
        END
        AntennaDiffArea 0.363 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.810 0.960 1.870 1.220 ;
        RECT  1.750 0.960 1.810 1.375 ;
        RECT  1.470 1.030 1.750 1.375 ;
        END
        AntennaGateArea 0.077 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.715 0.535 1.895 ;
        END
        AntennaGateArea 0.117 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.535 -0.210 7.000 0.210 ;
        RECT  6.365 -0.210 6.535 0.285 ;
        RECT  5.810 -0.210 6.365 0.210 ;
        RECT  5.580 -0.210 5.810 0.850 ;
        RECT  3.970 -0.210 5.580 0.210 ;
        RECT  3.450 -0.210 3.970 0.285 ;
        RECT  2.440 -0.210 3.450 0.210 ;
        RECT  2.180 -0.210 2.440 0.285 ;
        RECT  1.750 -0.210 2.180 0.210 ;
        RECT  1.490 -0.210 1.750 0.285 ;
        RECT  0.660 -0.210 1.490 0.210 ;
        RECT  0.400 -0.210 0.660 0.870 ;
        RECT  0.000 -0.210 0.400 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.535 2.310 7.000 2.730 ;
        RECT  6.365 2.260 6.535 2.730 ;
        RECT  5.735 2.310 6.365 2.730 ;
        RECT  5.565 2.260 5.735 2.730 ;
        RECT  3.965 2.310 5.565 2.730 ;
        RECT  3.445 2.220 3.965 2.730 ;
        RECT  2.165 2.310 3.445 2.730 ;
        RECT  1.735 2.175 2.165 2.730 ;
        RECT  0.610 2.310 1.735 2.730 ;
        RECT  0.350 2.015 0.610 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.610 1.020 6.670 1.280 ;
        RECT  6.490 1.020 6.610 2.140 ;
        RECT  6.180 2.020 6.490 2.140 ;
        RECT  6.185 0.635 6.255 0.805 ;
        RECT  6.185 1.460 6.230 1.720 ;
        RECT  6.065 0.635 6.185 1.720 ;
        RECT  5.920 2.020 6.180 2.190 ;
        RECT  5.630 1.005 6.065 1.265 ;
        RECT  5.695 2.020 5.920 2.140 ;
        RECT  5.575 1.530 5.695 2.140 ;
        RECT  5.160 1.530 5.575 1.650 ;
        RECT  5.400 1.150 5.460 1.410 ;
        RECT  5.280 0.405 5.400 1.410 ;
        RECT  4.550 0.405 5.280 0.525 ;
        RECT  5.040 0.660 5.160 1.650 ;
        RECT  4.840 0.660 5.040 0.780 ;
        RECT  4.680 1.345 4.840 1.840 ;
        RECT  4.545 1.960 4.715 2.145 ;
        RECT  4.410 0.660 4.680 1.840 ;
        RECT  4.290 0.375 4.550 0.525 ;
        RECT  2.800 1.960 4.545 2.080 ;
        RECT  4.160 0.660 4.410 0.780 ;
        RECT  2.660 1.720 4.410 1.840 ;
        RECT  3.595 0.405 4.290 0.525 ;
        RECT  4.145 0.940 4.190 1.200 ;
        RECT  4.025 0.940 4.145 1.595 ;
        RECT  3.305 1.475 4.025 1.595 ;
        RECT  3.475 0.405 3.595 1.355 ;
        RECT  2.830 0.405 3.475 0.525 ;
        RECT  3.425 1.185 3.475 1.355 ;
        RECT  3.185 0.730 3.305 1.595 ;
        RECT  2.980 0.730 3.185 0.850 ;
        RECT  2.780 1.475 3.185 1.595 ;
        RECT  2.940 0.990 3.060 1.250 ;
        RECT  2.720 0.660 2.980 0.850 ;
        RECT  2.600 0.990 2.940 1.110 ;
        RECT  2.570 0.350 2.830 0.525 ;
        RECT  2.540 1.960 2.800 2.150 ;
        RECT  2.540 1.470 2.660 1.840 ;
        RECT  2.480 0.675 2.600 1.110 ;
        RECT  0.950 0.405 2.570 0.525 ;
        RECT  2.360 1.470 2.540 1.590 ;
        RECT  2.420 1.960 2.540 2.080 ;
        RECT  2.110 0.675 2.480 0.795 ;
        RECT  2.300 1.720 2.420 2.080 ;
        RECT  2.240 1.035 2.360 1.590 ;
        RECT  1.190 1.720 2.300 1.840 ;
        RECT  1.990 0.675 2.110 1.600 ;
        RECT  1.830 0.675 1.990 0.820 ;
        RECT  1.930 1.340 1.990 1.600 ;
        RECT  1.100 1.990 1.360 2.170 ;
        RECT  1.190 0.675 1.325 0.845 ;
        RECT  1.070 0.675 1.190 1.840 ;
        RECT  0.920 1.990 1.100 2.110 ;
        RECT  1.040 1.470 1.070 1.730 ;
        RECT  0.920 0.405 0.950 0.920 ;
        RECT  0.800 0.405 0.920 2.110 ;
        RECT  0.740 1.850 0.800 2.110 ;
        RECT  0.255 1.020 0.680 1.280 ;
        RECT  0.135 0.680 0.255 1.555 ;
        RECT  0.110 0.680 0.135 0.940 ;
        RECT  0.085 1.385 0.135 1.555 ;
    END
END DFFHQX2AD
MACRO DFFHQX4AD
    CLASS CORE ;
    FOREIGN DFFHQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.940 1.005 8.050 1.515 ;
        RECT  7.810 0.410 7.940 2.005 ;
        END
        AntennaDiffArea 0.41 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.080 2.505 1.375 ;
        END
        AntennaGateArea 0.108 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.050 1.510 1.220 ;
        RECT  1.075 0.865 1.450 1.220 ;
        END
        AntennaGateArea 0.197 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.315 -0.210 8.400 0.210 ;
        RECT  8.145 -0.210 8.315 0.865 ;
        RECT  7.620 -0.210 8.145 0.210 ;
        RECT  7.360 -0.210 7.620 0.300 ;
        RECT  6.475 -0.210 7.360 0.210 ;
        RECT  6.305 -0.210 6.475 0.255 ;
        RECT  4.945 -0.210 6.305 0.210 ;
        RECT  4.685 -0.210 4.945 0.260 ;
        RECT  3.070 -0.210 4.685 0.210 ;
        RECT  2.810 -0.210 3.070 0.260 ;
        RECT  1.380 -0.210 2.810 0.210 ;
        RECT  1.120 -0.210 1.380 0.260 ;
        RECT  0.230 -0.210 1.120 0.210 ;
        RECT  0.110 -0.210 0.230 0.860 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.290 2.310 8.400 2.730 ;
        RECT  8.170 1.600 8.290 2.730 ;
        RECT  7.575 2.310 8.170 2.730 ;
        RECT  7.405 2.265 7.575 2.730 ;
        RECT  6.660 2.310 7.405 2.730 ;
        RECT  6.400 2.110 6.660 2.730 ;
        RECT  5.090 2.310 6.400 2.730 ;
        RECT  4.920 2.265 5.090 2.730 ;
        RECT  4.165 2.310 4.920 2.730 ;
        RECT  3.995 2.265 4.165 2.730 ;
        RECT  2.925 2.310 3.995 2.730 ;
        RECT  2.755 2.265 2.925 2.730 ;
        RECT  1.580 2.310 2.755 2.730 ;
        RECT  1.320 2.190 1.580 2.730 ;
        RECT  0.975 2.310 1.320 2.730 ;
        RECT  0.805 1.885 0.975 2.730 ;
        RECT  0.230 2.310 0.805 2.730 ;
        RECT  0.110 1.580 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.400 2.520 ;
        LAYER M1 ;
        RECT  7.570 0.485 7.690 1.980 ;
        RECT  7.150 0.485 7.570 0.605 ;
        RECT  7.310 1.860 7.570 1.980 ;
        RECT  7.050 1.860 7.310 2.070 ;
        RECT  7.115 0.760 7.285 1.740 ;
        RECT  6.890 0.330 7.150 0.605 ;
        RECT  6.620 0.760 7.115 0.880 ;
        RECT  6.590 1.620 7.115 1.740 ;
        RECT  6.450 1.860 7.050 1.980 ;
        RECT  6.380 1.290 6.995 1.410 ;
        RECT  6.500 0.570 6.620 0.880 ;
        RECT  6.330 1.530 6.450 1.980 ;
        RECT  6.260 0.380 6.380 1.410 ;
        RECT  5.875 1.530 6.330 1.650 ;
        RECT  5.550 0.380 6.260 0.500 ;
        RECT  6.090 1.770 6.210 2.030 ;
        RECT  5.360 0.620 6.120 0.740 ;
        RECT  5.515 1.770 6.090 1.895 ;
        RECT  5.845 1.480 5.875 1.650 ;
        RECT  5.705 0.865 5.845 1.650 ;
        RECT  5.670 2.070 5.730 2.190 ;
        RECT  5.480 0.865 5.705 0.985 ;
        RECT  5.470 2.020 5.670 2.190 ;
        RECT  5.290 0.330 5.550 0.500 ;
        RECT  5.360 1.690 5.515 1.895 ;
        RECT  3.380 2.020 5.470 2.140 ;
        RECT  5.240 0.620 5.360 1.895 ;
        RECT  4.480 0.380 5.290 0.500 ;
        RECT  5.080 0.670 5.240 0.790 ;
        RECT  3.000 1.770 5.240 1.895 ;
        RECT  4.785 0.975 5.120 1.235 ;
        RECT  4.665 0.880 4.785 1.650 ;
        RECT  4.360 0.880 4.665 1.000 ;
        RECT  3.295 1.530 4.665 1.650 ;
        RECT  4.410 1.150 4.530 1.410 ;
        RECT  4.220 0.330 4.480 0.500 ;
        RECT  3.255 1.260 4.410 1.410 ;
        RECT  4.240 0.620 4.360 1.000 ;
        RECT  3.580 0.620 4.240 0.740 ;
        RECT  0.615 0.380 4.220 0.500 ;
        RECT  3.120 2.020 3.380 2.190 ;
        RECT  3.135 0.620 3.255 1.410 ;
        RECT  2.760 0.620 3.135 0.740 ;
        RECT  2.760 2.020 3.120 2.140 ;
        RECT  2.880 1.150 3.000 1.895 ;
        RECT  2.640 0.620 2.760 1.650 ;
        RECT  2.640 1.780 2.760 2.140 ;
        RECT  2.330 0.620 2.640 0.740 ;
        RECT  2.330 1.530 2.640 1.650 ;
        RECT  2.165 1.780 2.640 1.900 ;
        RECT  2.140 2.020 2.400 2.190 ;
        RECT  1.995 1.690 2.165 1.900 ;
        RECT  1.820 2.020 2.140 2.140 ;
        RECT  1.750 1.690 1.995 1.810 ;
        RECT  1.700 1.930 1.820 2.140 ;
        RECT  1.630 0.680 1.750 1.810 ;
        RECT  1.260 1.930 1.700 2.050 ;
        RECT  1.570 0.680 1.630 0.940 ;
        RECT  0.955 1.400 1.290 1.520 ;
        RECT  1.140 1.640 1.260 2.050 ;
        RECT  0.615 1.640 1.140 1.760 ;
        RECT  0.835 0.680 0.955 1.520 ;
        RECT  0.785 0.680 0.835 1.260 ;
        RECT  0.620 1.000 0.785 1.260 ;
        RECT  0.475 0.380 0.615 0.810 ;
        RECT  0.475 1.610 0.615 2.040 ;
        RECT  0.445 0.380 0.475 2.040 ;
        RECT  0.350 0.640 0.445 2.040 ;
    END
END DFFHQX4AD
MACRO DFFHQX8AD
    CLASS CORE ;
    FOREIGN DFFHQX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.370 0.410 13.570 2.005 ;
        RECT  12.835 1.005 13.370 1.515 ;
        RECT  12.665 0.410 12.835 2.005 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.570 1.065 3.850 1.235 ;
        RECT  3.430 1.065 3.570 1.375 ;
        END
        AntennaGateArea 0.219 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.065 1.770 1.235 ;
        RECT  1.340 0.865 1.720 1.235 ;
        END
        AntennaGateArea 0.353 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.915 -0.210 14.000 0.210 ;
        RECT  13.745 -0.210 13.915 0.865 ;
        RECT  13.195 -0.210 13.745 0.210 ;
        RECT  13.025 -0.210 13.195 0.865 ;
        RECT  12.405 -0.210 13.025 0.210 ;
        RECT  12.235 -0.210 12.405 0.260 ;
        RECT  11.850 -0.210 12.235 0.210 ;
        RECT  11.680 -0.210 11.850 0.260 ;
        RECT  8.800 -0.210 11.680 0.210 ;
        RECT  8.630 -0.210 8.800 0.260 ;
        RECT  8.040 -0.210 8.630 0.210 ;
        RECT  7.870 -0.210 8.040 0.260 ;
        RECT  7.280 -0.210 7.870 0.210 ;
        RECT  7.110 -0.210 7.280 0.260 ;
        RECT  5.995 -0.210 7.110 0.210 ;
        RECT  5.735 -0.210 5.995 0.430 ;
        RECT  4.575 -0.210 5.735 0.210 ;
        RECT  4.405 -0.210 4.575 0.260 ;
        RECT  1.625 -0.210 4.405 0.210 ;
        RECT  1.455 -0.210 1.625 0.260 ;
        RECT  0.590 -0.210 1.455 0.210 ;
        RECT  0.470 -0.210 0.590 0.860 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.915 2.310 14.000 2.730 ;
        RECT  13.745 1.645 13.915 2.730 ;
        RECT  13.195 2.310 13.745 2.730 ;
        RECT  13.025 1.725 13.195 2.730 ;
        RECT  12.405 2.310 13.025 2.730 ;
        RECT  12.235 2.260 12.405 2.730 ;
        RECT  11.990 2.310 12.235 2.730 ;
        RECT  11.820 2.260 11.990 2.730 ;
        RECT  8.610 2.310 11.820 2.730 ;
        RECT  8.440 2.220 8.610 2.730 ;
        RECT  7.850 2.310 8.440 2.730 ;
        RECT  7.680 2.220 7.850 2.730 ;
        RECT  7.115 2.310 7.680 2.730 ;
        RECT  6.945 2.220 7.115 2.730 ;
        RECT  5.695 2.310 6.945 2.730 ;
        RECT  5.525 2.220 5.695 2.730 ;
        RECT  4.350 2.310 5.525 2.730 ;
        RECT  4.180 2.220 4.350 2.730 ;
        RECT  3.655 2.310 4.180 2.730 ;
        RECT  3.395 2.035 3.655 2.730 ;
        RECT  2.030 2.310 3.395 2.730 ;
        RECT  1.770 2.190 2.030 2.730 ;
        RECT  1.380 2.310 1.770 2.730 ;
        RECT  1.120 2.040 1.380 2.730 ;
        RECT  0.590 2.310 1.120 2.730 ;
        RECT  0.470 1.575 0.590 2.730 ;
        RECT  0.000 2.310 0.470 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 14.000 2.520 ;
        LAYER M1 ;
        RECT  12.410 1.060 12.530 2.140 ;
        RECT  12.360 1.060 12.410 1.230 ;
        RECT  11.490 2.020 12.410 2.140 ;
        RECT  12.090 0.760 12.210 1.590 ;
        RECT  11.950 0.760 12.090 1.165 ;
        RECT  12.020 1.330 12.090 1.590 ;
        RECT  11.690 0.995 11.950 1.165 ;
        RECT  11.450 0.380 11.570 1.725 ;
        RECT  11.370 1.845 11.490 2.140 ;
        RECT  9.090 0.380 11.450 0.500 ;
        RECT  11.290 1.845 11.370 1.965 ;
        RECT  11.170 0.640 11.290 1.965 ;
        RECT  11.075 0.640 11.170 0.985 ;
        RECT  9.515 1.505 11.170 1.625 ;
        RECT  9.500 0.865 11.075 0.985 ;
        RECT  8.360 0.620 10.925 0.740 ;
        RECT  9.465 1.785 10.860 1.905 ;
        RECT  9.365 1.740 9.465 1.905 ;
        RECT  8.360 1.740 9.365 1.860 ;
        RECT  8.965 1.980 9.225 2.145 ;
        RECT  8.920 0.330 9.090 0.500 ;
        RECT  4.895 1.980 8.965 2.100 ;
        RECT  6.240 0.380 8.920 0.500 ;
        RECT  8.240 0.620 8.360 1.860 ;
        RECT  7.445 0.620 8.240 0.740 ;
        RECT  7.515 1.740 8.240 1.860 ;
        RECT  6.840 0.950 8.105 1.070 ;
        RECT  7.255 1.400 7.515 1.860 ;
        RECT  7.040 1.660 7.255 1.860 ;
        RECT  4.495 1.740 7.040 1.860 ;
        RECT  6.720 0.690 6.840 1.620 ;
        RECT  6.525 0.690 6.720 0.910 ;
        RECT  4.850 1.500 6.720 1.620 ;
        RECT  5.190 1.030 6.600 1.190 ;
        RECT  5.265 0.790 6.525 0.910 ;
        RECT  6.120 0.380 6.240 0.670 ;
        RECT  5.575 0.550 6.120 0.670 ;
        RECT  5.455 0.380 5.575 0.670 ;
        RECT  1.020 0.380 5.455 0.500 ;
        RECT  5.005 0.700 5.265 0.910 ;
        RECT  5.070 1.030 5.190 1.290 ;
        RECT  4.170 1.030 5.070 1.150 ;
        RECT  4.635 1.980 4.895 2.190 ;
        RECT  4.255 1.980 4.635 2.100 ;
        RECT  4.375 1.300 4.495 1.860 ;
        RECT  4.135 1.740 4.255 2.100 ;
        RECT  4.050 0.630 4.170 1.620 ;
        RECT  2.965 1.740 4.135 1.860 ;
        RECT  3.755 1.500 4.050 1.620 ;
        RECT  2.445 1.690 2.965 1.860 ;
        RECT  2.590 1.980 2.850 2.190 ;
        RECT  2.270 1.980 2.590 2.100 ;
        RECT  2.050 1.690 2.445 1.810 ;
        RECT  2.150 1.930 2.270 2.100 ;
        RECT  1.620 1.930 2.150 2.050 ;
        RECT  1.930 0.670 2.050 1.810 ;
        RECT  1.860 0.670 1.930 0.930 ;
        RECT  1.220 1.500 1.650 1.660 ;
        RECT  1.500 1.800 1.620 2.050 ;
        RECT  0.975 1.800 1.500 1.920 ;
        RECT  1.100 0.690 1.220 1.660 ;
        RECT  0.980 1.000 1.100 1.260 ;
        RECT  0.835 0.380 1.020 0.550 ;
        RECT  0.835 1.620 0.975 2.050 ;
        RECT  0.710 0.380 0.835 2.050 ;
        RECT  0.230 1.145 0.710 1.265 ;
        RECT  0.110 0.510 0.230 2.095 ;
    END
END DFFHQX8AD
MACRO DFFHX1AD
    CLASS CORE ;
    FOREIGN DFFHX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.040 0.655 7.210 1.600 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.370 1.375 6.425 1.545 ;
        RECT  6.370 0.645 6.400 0.905 ;
        RECT  6.230 0.645 6.370 1.545 ;
        END
        AntennaDiffArea 0.213 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.000 1.890 1.260 ;
        RECT  1.610 1.100 1.770 1.260 ;
        RECT  1.470 1.100 1.610 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.170 1.715 0.535 1.890 ;
        END
        AntennaGateArea 0.114 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.815 -0.210 7.280 0.210 ;
        RECT  6.645 -0.210 6.815 0.870 ;
        RECT  5.775 -0.210 6.645 0.210 ;
        RECT  5.515 -0.210 5.775 0.370 ;
        RECT  3.930 -0.210 5.515 0.210 ;
        RECT  3.670 -0.210 3.930 0.300 ;
        RECT  2.560 -0.210 3.670 0.210 ;
        RECT  2.300 -0.210 2.560 0.300 ;
        RECT  1.765 -0.210 2.300 0.210 ;
        RECT  1.505 -0.210 1.765 0.300 ;
        RECT  0.600 -0.210 1.505 0.210 ;
        RECT  0.600 0.750 0.670 0.870 ;
        RECT  0.480 -0.210 0.600 0.870 ;
        RECT  0.000 -0.210 0.480 0.210 ;
        RECT  0.410 0.750 0.480 0.870 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.805 2.310 7.280 2.730 ;
        RECT  6.805 2.030 6.850 2.150 ;
        RECT  6.635 1.990 6.805 2.730 ;
        RECT  6.590 2.030 6.635 2.150 ;
        RECT  5.740 2.310 6.635 2.730 ;
        RECT  5.480 2.180 5.740 2.730 ;
        RECT  4.165 2.310 5.480 2.730 ;
        RECT  3.645 2.220 4.165 2.730 ;
        RECT  2.105 2.310 3.645 2.730 ;
        RECT  1.675 1.950 2.105 2.730 ;
        RECT  0.600 2.310 1.675 2.730 ;
        RECT  0.340 2.010 0.600 2.730 ;
        RECT  0.000 2.310 0.340 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.280 2.520 ;
        LAYER M1 ;
        RECT  6.800 1.020 6.920 1.785 ;
        RECT  6.050 1.665 6.800 1.785 ;
        RECT  5.930 0.550 6.050 1.785 ;
        RECT  5.810 1.905 6.000 2.025 ;
        RECT  5.570 0.860 5.930 0.980 ;
        RECT  5.690 1.480 5.810 2.025 ;
        RECT  4.910 1.480 5.690 1.600 ;
        RECT  5.450 0.860 5.570 1.120 ;
        RECT  5.150 1.100 5.180 1.360 ;
        RECT  4.900 1.960 5.160 2.170 ;
        RECT  5.070 0.380 5.150 1.360 ;
        RECT  5.030 0.330 5.070 1.360 ;
        RECT  4.810 0.330 5.030 0.500 ;
        RECT  4.790 0.620 4.910 1.820 ;
        RECT  2.345 1.960 4.900 2.080 ;
        RECT  4.140 0.380 4.810 0.500 ;
        RECT  4.650 0.620 4.790 0.740 ;
        RECT  4.505 1.400 4.555 1.830 ;
        RECT  4.385 0.620 4.505 1.830 ;
        RECT  4.230 0.620 4.385 0.740 ;
        RECT  2.600 1.710 4.385 1.830 ;
        RECT  4.145 0.880 4.265 1.140 ;
        RECT  4.030 1.020 4.145 1.140 ;
        RECT  4.020 0.380 4.140 0.540 ;
        RECT  3.910 1.020 4.030 1.590 ;
        RECT  3.690 0.420 4.020 0.540 ;
        RECT  3.450 1.470 3.910 1.590 ;
        RECT  3.570 0.420 3.690 1.350 ;
        RECT  3.040 0.420 3.570 0.540 ;
        RECT  3.330 0.730 3.450 1.590 ;
        RECT  3.210 0.730 3.330 0.850 ;
        RECT  2.950 1.410 3.330 1.590 ;
        RECT  2.950 0.670 3.210 0.850 ;
        RECT  3.090 0.990 3.210 1.250 ;
        RECT  2.830 0.990 3.090 1.110 ;
        RECT  2.780 0.360 3.040 0.540 ;
        RECT  2.710 0.680 2.830 1.110 ;
        RECT  0.960 0.420 2.780 0.540 ;
        RECT  2.130 0.680 2.710 0.800 ;
        RECT  2.570 1.470 2.600 1.830 ;
        RECT  2.480 0.970 2.570 1.830 ;
        RECT  2.420 0.970 2.480 1.590 ;
        RECT  2.225 1.710 2.345 2.080 ;
        RECT  1.270 1.710 2.225 1.830 ;
        RECT  2.010 0.680 2.130 1.590 ;
        RECT  1.850 0.680 2.010 0.860 ;
        RECT  1.120 1.950 1.380 2.170 ;
        RECT  1.270 0.675 1.335 0.845 ;
        RECT  1.150 0.675 1.270 1.830 ;
        RECT  1.060 1.410 1.150 1.670 ;
        RECT  0.990 1.950 1.120 2.070 ;
        RECT  0.930 1.845 0.990 2.070 ;
        RECT  0.930 0.420 0.960 0.920 ;
        RECT  0.810 0.420 0.930 2.070 ;
        RECT  0.775 1.845 0.810 2.070 ;
        RECT  0.730 1.845 0.775 1.965 ;
        RECT  0.570 0.990 0.690 1.250 ;
        RECT  0.265 1.060 0.570 1.180 ;
        RECT  0.240 0.815 0.265 1.595 ;
        RECT  0.145 0.680 0.240 1.595 ;
        RECT  0.120 0.680 0.145 0.940 ;
        RECT  0.120 1.335 0.145 1.595 ;
    END
END DFFHX1AD
MACRO DFFHX2AD
    CLASS CORE ;
    FOREIGN DFFHX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.790 0.405 6.930 1.900 ;
        RECT  6.760 0.405 6.790 0.525 ;
        RECT  6.500 1.780 6.790 1.900 ;
        RECT  6.500 0.330 6.760 0.525 ;
        END
        AntennaDiffArea 0.126 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 0.685 7.490 1.580 ;
        RECT  7.350 0.355 7.450 2.170 ;
        RECT  7.290 0.355 7.350 0.875 ;
        RECT  7.290 1.390 7.350 2.170 ;
        END
        AntennaDiffArea 0.363 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.810 0.960 1.870 1.220 ;
        RECT  1.750 0.960 1.810 1.375 ;
        RECT  1.470 1.030 1.750 1.375 ;
        END
        AntennaGateArea 0.049 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.715 0.535 1.895 ;
        END
        AntennaGateArea 0.125 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.095 -0.210 7.560 0.210 ;
        RECT  6.925 -0.210 7.095 0.285 ;
        RECT  6.240 -0.210 6.925 0.210 ;
        RECT  6.070 -0.210 6.240 0.815 ;
        RECT  4.760 -0.210 6.070 0.210 ;
        RECT  4.500 -0.210 4.760 0.285 ;
        RECT  3.970 -0.210 4.500 0.210 ;
        RECT  3.450 -0.210 3.970 0.285 ;
        RECT  2.440 -0.210 3.450 0.210 ;
        RECT  2.180 -0.210 2.440 0.285 ;
        RECT  1.750 -0.210 2.180 0.210 ;
        RECT  1.490 -0.210 1.750 0.285 ;
        RECT  0.660 -0.210 1.490 0.210 ;
        RECT  0.400 -0.210 0.660 0.870 ;
        RECT  0.000 -0.210 0.400 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.095 2.310 7.560 2.730 ;
        RECT  6.925 2.260 7.095 2.730 ;
        RECT  6.095 2.310 6.925 2.730 ;
        RECT  5.925 2.260 6.095 2.730 ;
        RECT  4.750 2.310 5.925 2.730 ;
        RECT  4.490 2.220 4.750 2.730 ;
        RECT  4.230 2.310 4.490 2.730 ;
        RECT  3.970 2.220 4.230 2.730 ;
        RECT  3.705 2.310 3.970 2.730 ;
        RECT  3.445 2.220 3.705 2.730 ;
        RECT  2.165 2.310 3.445 2.730 ;
        RECT  1.735 1.960 2.165 2.730 ;
        RECT  0.610 2.310 1.735 2.730 ;
        RECT  0.350 2.015 0.610 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  7.170 1.020 7.230 1.280 ;
        RECT  7.050 1.020 7.170 2.140 ;
        RECT  6.540 2.020 7.050 2.140 ;
        RECT  6.565 1.290 6.630 1.550 ;
        RECT  6.565 0.645 6.615 0.815 ;
        RECT  6.445 0.645 6.565 1.550 ;
        RECT  6.280 2.020 6.540 2.190 ;
        RECT  6.010 1.005 6.445 1.265 ;
        RECT  5.790 2.020 6.280 2.140 ;
        RECT  5.730 0.405 5.850 1.410 ;
        RECT  5.580 1.960 5.790 2.140 ;
        RECT  5.000 0.405 5.730 0.525 ;
        RECT  5.700 1.150 5.730 1.410 ;
        RECT  5.580 0.645 5.605 0.815 ;
        RECT  5.460 0.645 5.580 2.140 ;
        RECT  5.435 0.645 5.460 0.815 ;
        RECT  5.315 1.460 5.340 1.980 ;
        RECT  5.220 0.710 5.315 1.980 ;
        RECT  5.195 0.710 5.220 1.895 ;
        RECT  4.435 0.710 5.195 0.830 ;
        RECT  4.930 1.150 5.050 2.080 ;
        RECT  4.720 0.405 5.000 0.570 ;
        RECT  2.800 1.960 4.930 2.080 ;
        RECT  3.595 0.405 4.720 0.525 ;
        RECT  4.315 0.680 4.435 1.840 ;
        RECT  4.110 0.680 4.315 0.800 ;
        RECT  4.265 1.345 4.315 1.840 ;
        RECT  2.660 1.720 4.265 1.840 ;
        RECT  4.145 0.940 4.190 1.200 ;
        RECT  4.025 0.940 4.145 1.595 ;
        RECT  3.305 1.475 4.025 1.595 ;
        RECT  3.475 0.405 3.595 1.355 ;
        RECT  2.830 0.405 3.475 0.525 ;
        RECT  3.425 1.185 3.475 1.355 ;
        RECT  3.185 0.730 3.305 1.595 ;
        RECT  2.980 0.730 3.185 0.850 ;
        RECT  2.780 1.475 3.185 1.595 ;
        RECT  2.940 0.990 3.060 1.250 ;
        RECT  2.720 0.680 2.980 0.850 ;
        RECT  2.600 0.990 2.940 1.110 ;
        RECT  2.570 0.370 2.830 0.525 ;
        RECT  2.540 1.960 2.800 2.150 ;
        RECT  2.540 1.470 2.660 1.840 ;
        RECT  2.480 0.675 2.600 1.110 ;
        RECT  0.950 0.405 2.570 0.525 ;
        RECT  2.360 1.470 2.540 1.590 ;
        RECT  2.420 1.960 2.540 2.080 ;
        RECT  2.110 0.675 2.480 0.795 ;
        RECT  2.300 1.720 2.420 2.080 ;
        RECT  2.240 1.035 2.360 1.590 ;
        RECT  1.190 1.720 2.300 1.840 ;
        RECT  1.990 0.675 2.110 1.600 ;
        RECT  1.830 0.675 1.990 0.820 ;
        RECT  1.930 1.340 1.990 1.600 ;
        RECT  1.100 1.990 1.360 2.170 ;
        RECT  1.190 0.675 1.325 0.845 ;
        RECT  1.070 0.675 1.190 1.840 ;
        RECT  0.920 1.990 1.100 2.110 ;
        RECT  1.040 1.470 1.070 1.730 ;
        RECT  0.920 0.405 0.950 0.920 ;
        RECT  0.800 0.405 0.920 2.110 ;
        RECT  0.740 1.850 0.800 2.110 ;
        RECT  0.255 1.020 0.680 1.280 ;
        RECT  0.135 0.680 0.255 1.555 ;
        RECT  0.110 0.680 0.135 0.940 ;
        RECT  0.085 1.385 0.135 1.555 ;
    END
END DFFHX2AD
MACRO DFFHX4AD
    CLASS CORE ;
    FOREIGN DFFHX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.555 1.750 7.955 1.900 ;
        RECT  7.555 0.760 7.770 0.890 ;
        RECT  7.425 0.760 7.555 1.900 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.500 1.005 8.610 1.515 ;
        RECT  8.370 0.410 8.500 2.005 ;
        END
        AntennaDiffArea 0.41 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.130 2.510 1.390 ;
        END
        AntennaGateArea 0.076 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.050 1.510 1.220 ;
        RECT  1.075 0.865 1.450 1.220 ;
        END
        AntennaGateArea 0.197 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.875 -0.210 8.960 0.210 ;
        RECT  8.705 -0.210 8.875 0.865 ;
        RECT  8.180 -0.210 8.705 0.210 ;
        RECT  7.920 -0.210 8.180 0.300 ;
        RECT  7.380 -0.210 7.920 0.210 ;
        RECT  7.120 -0.210 7.380 0.300 ;
        RECT  6.530 -0.210 7.120 0.210 ;
        RECT  6.360 -0.210 6.530 0.260 ;
        RECT  4.990 -0.210 6.360 0.210 ;
        RECT  4.730 -0.210 4.990 0.260 ;
        RECT  3.080 -0.210 4.730 0.210 ;
        RECT  2.820 -0.210 3.080 0.260 ;
        RECT  1.380 -0.210 2.820 0.210 ;
        RECT  1.120 -0.210 1.380 0.260 ;
        RECT  0.230 -0.210 1.120 0.210 ;
        RECT  0.110 -0.210 0.230 0.860 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.850 2.310 8.960 2.730 ;
        RECT  8.730 1.600 8.850 2.730 ;
        RECT  8.135 2.310 8.730 2.730 ;
        RECT  7.965 2.265 8.135 2.730 ;
        RECT  7.445 2.310 7.965 2.730 ;
        RECT  7.275 2.265 7.445 2.730 ;
        RECT  6.695 2.310 7.275 2.730 ;
        RECT  6.435 2.220 6.695 2.730 ;
        RECT  5.055 2.310 6.435 2.730 ;
        RECT  4.885 2.265 5.055 2.730 ;
        RECT  4.155 2.310 4.885 2.730 ;
        RECT  3.985 2.265 4.155 2.730 ;
        RECT  2.915 2.310 3.985 2.730 ;
        RECT  2.745 2.265 2.915 2.730 ;
        RECT  1.580 2.310 2.745 2.730 ;
        RECT  1.320 2.190 1.580 2.730 ;
        RECT  0.975 2.310 1.320 2.730 ;
        RECT  0.805 1.885 0.975 2.730 ;
        RECT  0.230 2.310 0.805 2.730 ;
        RECT  0.110 1.580 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.960 2.520 ;
        LAYER M1 ;
        RECT  8.130 0.990 8.250 2.140 ;
        RECT  7.230 2.020 8.130 2.140 ;
        RECT  7.890 0.420 8.010 1.545 ;
        RECT  7.290 0.420 7.890 0.540 ;
        RECT  7.675 1.375 7.890 1.545 ;
        RECT  7.170 0.420 7.290 1.230 ;
        RECT  7.110 1.750 7.230 2.140 ;
        RECT  7.140 0.970 7.170 1.230 ;
        RECT  6.770 1.750 7.110 1.870 ;
        RECT  6.890 0.380 7.010 1.620 ;
        RECT  5.625 0.380 6.890 0.500 ;
        RECT  6.650 0.690 6.770 1.870 ;
        RECT  5.870 1.480 6.650 1.600 ;
        RECT  6.060 1.770 6.230 1.950 ;
        RECT  5.425 0.620 6.195 0.740 ;
        RECT  5.545 1.770 6.060 1.895 ;
        RECT  5.805 1.480 5.870 1.650 ;
        RECT  5.665 0.865 5.805 1.650 ;
        RECT  5.465 2.020 5.725 2.190 ;
        RECT  5.545 0.865 5.665 0.985 ;
        RECT  5.365 0.330 5.625 0.500 ;
        RECT  5.425 1.690 5.545 1.895 ;
        RECT  3.360 2.020 5.465 2.140 ;
        RECT  5.305 0.620 5.425 1.895 ;
        RECT  4.480 0.380 5.365 0.500 ;
        RECT  5.125 0.670 5.305 0.790 ;
        RECT  5.015 1.770 5.305 1.895 ;
        RECT  4.810 0.950 5.170 1.070 ;
        RECT  4.895 1.215 5.015 1.895 ;
        RECT  2.990 1.770 4.895 1.895 ;
        RECT  4.775 0.880 4.810 1.070 ;
        RECT  4.655 0.880 4.775 1.650 ;
        RECT  4.360 0.880 4.655 1.000 ;
        RECT  3.295 1.530 4.655 1.650 ;
        RECT  4.400 1.150 4.520 1.410 ;
        RECT  4.220 0.330 4.480 0.500 ;
        RECT  3.690 1.290 4.400 1.410 ;
        RECT  4.240 0.620 4.360 1.000 ;
        RECT  3.580 0.620 4.240 0.740 ;
        RECT  0.615 0.380 4.220 0.500 ;
        RECT  3.230 1.260 3.690 1.410 ;
        RECT  3.100 2.020 3.360 2.190 ;
        RECT  3.110 0.640 3.230 1.410 ;
        RECT  2.750 0.640 3.110 0.760 ;
        RECT  2.750 2.020 3.100 2.140 ;
        RECT  2.870 1.150 2.990 1.895 ;
        RECT  2.630 0.640 2.750 1.650 ;
        RECT  2.630 1.780 2.750 2.140 ;
        RECT  2.320 0.640 2.630 0.760 ;
        RECT  2.320 1.530 2.630 1.650 ;
        RECT  2.165 1.780 2.630 1.900 ;
        RECT  2.140 2.020 2.400 2.190 ;
        RECT  1.995 1.690 2.165 1.900 ;
        RECT  1.820 2.020 2.140 2.140 ;
        RECT  1.750 1.690 1.995 1.810 ;
        RECT  1.700 1.930 1.820 2.140 ;
        RECT  1.630 0.680 1.750 1.810 ;
        RECT  1.260 1.930 1.700 2.050 ;
        RECT  1.570 0.680 1.630 0.940 ;
        RECT  0.955 1.400 1.290 1.520 ;
        RECT  1.140 1.640 1.260 2.050 ;
        RECT  0.615 1.640 1.140 1.760 ;
        RECT  0.835 0.680 0.955 1.520 ;
        RECT  0.785 0.680 0.835 1.260 ;
        RECT  0.620 1.000 0.785 1.260 ;
        RECT  0.475 0.380 0.615 0.810 ;
        RECT  0.475 1.610 0.615 2.040 ;
        RECT  0.445 0.380 0.475 2.040 ;
        RECT  0.350 0.640 0.445 2.040 ;
    END
END DFFHX4AD
MACRO DFFHX8AD
    CLASS CORE ;
    FOREIGN DFFHX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.280 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.175 1.740 12.415 1.900 ;
        RECT  12.175 0.640 12.205 0.900 ;
        RECT  12.005 0.640 12.175 1.900 ;
        RECT  11.685 1.285 12.005 1.900 ;
        END
        AntennaDiffArea 0.124 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.650 0.410 13.850 2.005 ;
        RECT  13.115 1.005 13.650 1.515 ;
        RECT  12.945 0.410 13.115 2.005 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 1.065 3.820 1.375 ;
        END
        AntennaGateArea 0.139 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.065 1.770 1.235 ;
        RECT  1.340 0.865 1.720 1.235 ;
        END
        AntennaGateArea 0.353 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.195 -0.210 14.280 0.210 ;
        RECT  14.025 -0.210 14.195 0.865 ;
        RECT  13.475 -0.210 14.025 0.210 ;
        RECT  13.305 -0.210 13.475 0.865 ;
        RECT  12.730 -0.210 13.305 0.210 ;
        RECT  12.610 -0.210 12.730 0.720 ;
        RECT  11.850 -0.210 12.610 0.210 ;
        RECT  11.680 -0.210 11.850 0.260 ;
        RECT  8.800 -0.210 11.680 0.210 ;
        RECT  8.630 -0.210 8.800 0.260 ;
        RECT  8.040 -0.210 8.630 0.210 ;
        RECT  7.870 -0.210 8.040 0.260 ;
        RECT  7.280 -0.210 7.870 0.210 ;
        RECT  7.110 -0.210 7.280 0.260 ;
        RECT  5.900 -0.210 7.110 0.210 ;
        RECT  5.640 -0.210 5.900 0.430 ;
        RECT  4.490 -0.210 5.640 0.210 ;
        RECT  4.320 -0.210 4.490 0.260 ;
        RECT  1.625 -0.210 4.320 0.210 ;
        RECT  1.455 -0.210 1.625 0.260 ;
        RECT  0.590 -0.210 1.455 0.210 ;
        RECT  0.470 -0.210 0.590 0.860 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.195 2.310 14.280 2.730 ;
        RECT  14.025 1.645 14.195 2.730 ;
        RECT  13.475 2.310 14.025 2.730 ;
        RECT  13.305 1.725 13.475 2.730 ;
        RECT  12.685 2.310 13.305 2.730 ;
        RECT  12.515 2.260 12.685 2.730 ;
        RECT  11.990 2.310 12.515 2.730 ;
        RECT  11.820 2.260 11.990 2.730 ;
        RECT  8.610 2.310 11.820 2.730 ;
        RECT  8.440 2.220 8.610 2.730 ;
        RECT  7.850 2.310 8.440 2.730 ;
        RECT  7.680 2.220 7.850 2.730 ;
        RECT  7.115 2.310 7.680 2.730 ;
        RECT  6.945 2.220 7.115 2.730 ;
        RECT  5.640 2.310 6.945 2.730 ;
        RECT  5.470 2.220 5.640 2.730 ;
        RECT  4.305 2.310 5.470 2.730 ;
        RECT  4.135 2.220 4.305 2.730 ;
        RECT  3.650 2.310 4.135 2.730 ;
        RECT  3.390 2.035 3.650 2.730 ;
        RECT  2.030 2.310 3.390 2.730 ;
        RECT  1.770 2.190 2.030 2.730 ;
        RECT  1.380 2.310 1.770 2.730 ;
        RECT  1.120 2.040 1.380 2.730 ;
        RECT  0.590 2.310 1.120 2.730 ;
        RECT  0.470 1.575 0.590 2.730 ;
        RECT  0.000 2.310 0.470 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 14.280 2.520 ;
        LAYER M1 ;
        RECT  12.690 1.060 12.810 2.140 ;
        RECT  12.640 1.060 12.690 1.230 ;
        RECT  11.490 2.020 12.690 2.140 ;
        RECT  12.370 0.400 12.490 1.590 ;
        RECT  12.350 0.400 12.370 0.520 ;
        RECT  12.300 1.330 12.370 1.590 ;
        RECT  12.090 0.365 12.350 0.520 ;
        RECT  11.750 0.400 12.090 0.520 ;
        RECT  11.630 0.400 11.750 1.165 ;
        RECT  11.580 0.995 11.630 1.165 ;
        RECT  11.460 1.465 11.565 1.725 ;
        RECT  11.370 1.845 11.490 2.140 ;
        RECT  11.340 0.380 11.460 1.725 ;
        RECT  11.220 1.845 11.370 1.965 ;
        RECT  9.090 0.380 11.340 0.500 ;
        RECT  11.100 0.640 11.220 1.965 ;
        RECT  11.075 0.640 11.100 0.985 ;
        RECT  9.515 1.505 11.100 1.625 ;
        RECT  9.500 0.865 11.075 0.985 ;
        RECT  8.360 0.620 10.925 0.740 ;
        RECT  10.645 1.785 10.815 1.955 ;
        RECT  9.465 1.785 10.645 1.905 ;
        RECT  9.365 1.740 9.465 1.905 ;
        RECT  8.360 1.740 9.365 1.860 ;
        RECT  8.965 1.980 9.225 2.145 ;
        RECT  8.920 0.330 9.090 0.500 ;
        RECT  4.810 1.980 8.965 2.100 ;
        RECT  6.240 0.380 8.920 0.500 ;
        RECT  8.240 0.620 8.360 1.860 ;
        RECT  7.445 0.620 8.240 0.740 ;
        RECT  7.515 1.740 8.240 1.860 ;
        RECT  6.840 0.950 8.105 1.070 ;
        RECT  7.255 1.400 7.515 1.860 ;
        RECT  7.040 1.660 7.255 1.860 ;
        RECT  4.400 1.740 7.040 1.860 ;
        RECT  6.720 0.690 6.840 1.620 ;
        RECT  6.470 0.690 6.720 0.910 ;
        RECT  4.690 1.500 6.720 1.620 ;
        RECT  5.080 1.030 6.600 1.190 ;
        RECT  5.180 0.790 6.470 0.910 ;
        RECT  6.120 0.380 6.240 0.670 ;
        RECT  5.480 0.550 6.120 0.670 ;
        RECT  5.360 0.380 5.480 0.670 ;
        RECT  1.020 0.380 5.360 0.500 ;
        RECT  4.920 0.700 5.180 0.910 ;
        RECT  4.960 1.030 5.080 1.290 ;
        RECT  4.060 1.030 4.960 1.150 ;
        RECT  4.550 1.980 4.810 2.190 ;
        RECT  3.890 1.980 4.550 2.100 ;
        RECT  4.280 1.300 4.400 1.860 ;
        RECT  4.060 0.675 4.110 0.845 ;
        RECT  3.940 0.675 4.060 1.620 ;
        RECT  3.660 1.500 3.940 1.620 ;
        RECT  3.770 1.740 3.890 2.100 ;
        RECT  2.965 1.740 3.770 1.860 ;
        RECT  2.445 1.690 2.965 1.860 ;
        RECT  2.590 1.980 2.850 2.190 ;
        RECT  2.270 1.980 2.590 2.100 ;
        RECT  2.050 1.690 2.445 1.810 ;
        RECT  2.150 1.930 2.270 2.100 ;
        RECT  1.620 1.930 2.150 2.050 ;
        RECT  1.930 0.670 2.050 1.810 ;
        RECT  1.860 0.670 1.930 0.930 ;
        RECT  1.220 1.500 1.650 1.660 ;
        RECT  1.500 1.800 1.620 2.050 ;
        RECT  0.975 1.800 1.500 1.920 ;
        RECT  1.100 0.690 1.220 1.660 ;
        RECT  0.980 1.000 1.100 1.260 ;
        RECT  0.835 0.380 1.020 0.550 ;
        RECT  0.835 1.620 0.975 2.050 ;
        RECT  0.710 0.380 0.835 2.050 ;
        RECT  0.230 1.145 0.710 1.265 ;
        RECT  0.110 0.510 0.230 2.095 ;
    END
END DFFHX8AD
MACRO DFFNHX1AD
    CLASS CORE ;
    FOREIGN DFFNHX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.810 0.735 5.955 0.905 ;
        RECT  5.810 1.750 5.875 1.870 ;
        RECT  5.670 0.735 5.810 1.870 ;
        RECT  5.615 1.750 5.670 1.870 ;
        END
        AntennaDiffArea 0.139 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.875 1.145 6.930 1.375 ;
        RECT  6.750 0.610 6.875 1.925 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 0.910 2.215 1.205 ;
        END
        AntennaGateArea 0.061 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.175 1.045 1.330 1.375 ;
        RECT  1.095 1.045 1.175 1.305 ;
        END
        AntennaGateArea 0.118 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.565 -0.210 7.000 0.210 ;
        RECT  6.305 -0.210 6.565 0.310 ;
        RECT  5.615 -0.210 6.305 0.210 ;
        RECT  5.355 -0.210 5.615 0.285 ;
        RECT  4.125 -0.210 5.355 0.210 ;
        RECT  3.865 -0.210 4.125 0.300 ;
        RECT  2.420 -0.210 3.865 0.210 ;
        RECT  2.160 -0.210 2.420 0.300 ;
        RECT  1.325 -0.210 2.160 0.210 ;
        RECT  1.065 -0.210 1.325 0.430 ;
        RECT  0.285 -0.210 1.065 0.210 ;
        RECT  0.115 -0.210 0.285 0.875 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.565 2.310 7.000 2.730 ;
        RECT  6.305 1.925 6.565 2.730 ;
        RECT  5.495 2.310 6.305 2.730 ;
        RECT  5.235 2.230 5.495 2.730 ;
        RECT  4.015 2.310 5.235 2.730 ;
        RECT  3.755 2.220 4.015 2.730 ;
        RECT  2.765 2.310 3.755 2.730 ;
        RECT  2.505 2.220 2.765 2.730 ;
        RECT  1.335 2.310 2.505 2.730 ;
        RECT  1.075 1.965 1.335 2.730 ;
        RECT  0.285 2.310 1.075 2.730 ;
        RECT  0.115 1.540 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.500 1.050 6.550 1.220 ;
        RECT  6.380 1.050 6.500 1.785 ;
        RECT  6.125 1.665 6.380 1.785 ;
        RECT  6.095 0.405 6.215 1.545 ;
        RECT  6.005 1.665 6.125 2.110 ;
        RECT  5.550 0.405 6.095 0.525 ;
        RECT  5.965 1.375 6.095 1.545 ;
        RECT  4.980 1.990 6.005 2.110 ;
        RECT  5.430 0.405 5.550 1.580 ;
        RECT  5.015 0.420 5.135 1.600 ;
        RECT  4.825 0.420 5.015 0.540 ;
        RECT  4.775 1.480 5.015 1.600 ;
        RECT  4.860 1.780 4.980 2.110 ;
        RECT  4.715 0.690 4.875 1.050 ;
        RECT  4.655 1.780 4.860 1.900 ;
        RECT  4.565 0.330 4.825 0.540 ;
        RECT  4.655 0.930 4.715 1.050 ;
        RECT  4.535 0.930 4.655 1.900 ;
        RECT  4.410 0.690 4.585 0.810 ;
        RECT  3.645 0.420 4.565 0.540 ;
        RECT  4.350 2.070 4.555 2.190 ;
        RECT  4.290 0.690 4.410 1.860 ;
        RECT  4.230 1.980 4.350 2.190 ;
        RECT  4.075 0.690 4.290 0.810 ;
        RECT  4.190 1.570 4.290 1.860 ;
        RECT  3.245 1.980 4.230 2.100 ;
        RECT  2.855 1.740 4.190 1.860 ;
        RECT  3.605 1.190 4.170 1.310 ;
        RECT  3.815 0.690 4.075 0.980 ;
        RECT  3.525 0.380 3.645 0.540 ;
        RECT  3.485 0.660 3.605 1.620 ;
        RECT  3.240 0.380 3.525 0.500 ;
        RECT  3.405 0.660 3.485 0.780 ;
        RECT  3.115 1.500 3.485 1.620 ;
        RECT  3.255 0.620 3.405 0.780 ;
        RECT  3.235 1.065 3.355 1.330 ;
        RECT  2.845 0.620 3.255 0.740 ;
        RECT  2.985 1.980 3.245 2.140 ;
        RECT  2.980 0.330 3.240 0.500 ;
        RECT  2.475 1.065 3.235 1.185 ;
        RECT  2.190 1.980 2.985 2.100 ;
        RECT  2.740 0.380 2.980 0.500 ;
        RECT  2.735 1.360 2.855 1.860 ;
        RECT  2.620 0.380 2.740 0.540 ;
        RECT  2.595 1.360 2.735 1.480 ;
        RECT  1.655 0.420 2.620 0.540 ;
        RECT  2.375 0.660 2.475 1.570 ;
        RECT  2.355 0.660 2.375 1.810 ;
        RECT  1.815 0.660 2.355 0.780 ;
        RECT  2.255 1.450 2.355 1.810 ;
        RECT  2.115 1.690 2.255 1.810 ;
        RECT  2.070 1.980 2.190 2.140 ;
        RECT  1.845 2.020 2.070 2.140 ;
        RECT  1.775 1.380 1.895 1.900 ;
        RECT  1.650 2.020 1.845 2.190 ;
        RECT  1.655 1.380 1.775 1.500 ;
        RECT  1.535 0.420 1.655 1.500 ;
        RECT  1.530 1.725 1.650 2.190 ;
        RECT  0.645 1.725 1.530 1.845 ;
        RECT  0.975 1.425 1.000 1.595 ;
        RECT  0.855 0.680 0.975 1.595 ;
        RECT  0.830 1.020 0.855 1.595 ;
        RECT  0.755 1.020 0.830 1.280 ;
        RECT  0.620 1.540 0.645 1.970 ;
        RECT  0.500 0.660 0.620 1.970 ;
        RECT  0.475 1.540 0.500 1.970 ;
    END
END DFFNHX1AD
MACRO DFFNHX2AD
    CLASS CORE ;
    FOREIGN DFFNHX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.810 1.740 5.990 1.860 ;
        RECT  5.810 0.690 5.920 0.950 ;
        RECT  5.670 0.690 5.810 1.860 ;
        END
        AntennaDiffArea 0.133 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.875 0.735 6.930 1.625 ;
        RECT  6.790 0.400 6.875 2.145 ;
        RECT  6.705 0.400 6.790 0.830 ;
        RECT  6.705 1.455 6.790 2.145 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 0.910 2.215 1.225 ;
        END
        AntennaGateArea 0.087 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.175 1.045 1.330 1.375 ;
        RECT  1.095 1.045 1.175 1.305 ;
        END
        AntennaGateArea 0.127 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.515 -0.210 7.000 0.210 ;
        RECT  6.345 -0.210 6.515 0.555 ;
        RECT  5.610 -0.210 6.345 0.210 ;
        RECT  5.350 -0.210 5.610 0.300 ;
        RECT  4.160 -0.210 5.350 0.210 ;
        RECT  3.900 -0.210 4.160 0.290 ;
        RECT  2.370 -0.210 3.900 0.210 ;
        RECT  2.110 -0.210 2.370 0.290 ;
        RECT  1.325 -0.210 2.110 0.210 ;
        RECT  1.065 -0.210 1.325 0.365 ;
        RECT  0.285 -0.210 1.065 0.210 ;
        RECT  0.115 -0.210 0.285 0.875 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.520 2.310 7.000 2.730 ;
        RECT  6.350 1.885 6.520 2.730 ;
        RECT  5.610 2.310 6.350 2.730 ;
        RECT  5.350 2.220 5.610 2.730 ;
        RECT  4.115 2.310 5.350 2.730 ;
        RECT  3.855 2.230 4.115 2.730 ;
        RECT  2.685 2.310 3.855 2.730 ;
        RECT  2.425 2.230 2.685 2.730 ;
        RECT  1.335 2.310 2.425 2.730 ;
        RECT  1.075 1.965 1.335 2.730 ;
        RECT  0.285 2.310 1.075 2.730 ;
        RECT  0.115 1.480 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.440 1.045 6.560 1.760 ;
        RECT  6.355 1.045 6.440 1.215 ;
        RECT  6.230 1.640 6.440 1.760 ;
        RECT  6.160 1.400 6.250 1.520 ;
        RECT  6.110 1.640 6.230 2.100 ;
        RECT  6.040 0.385 6.160 1.520 ;
        RECT  5.305 1.980 6.110 2.100 ;
        RECT  5.985 0.385 6.040 0.555 ;
        RECT  5.990 1.400 6.040 1.520 ;
        RECT  5.410 0.435 5.985 0.555 ;
        RECT  5.290 0.435 5.410 1.525 ;
        RECT  5.185 1.670 5.305 2.100 ;
        RECT  4.665 1.670 5.185 1.790 ;
        RECT  5.025 0.330 5.145 1.510 ;
        RECT  4.785 1.980 5.045 2.190 ;
        RECT  4.885 0.330 5.025 0.500 ;
        RECT  4.875 1.390 5.025 1.510 ;
        RECT  4.855 0.645 4.905 0.815 ;
        RECT  4.415 0.380 4.885 0.500 ;
        RECT  4.735 0.645 4.855 1.080 ;
        RECT  3.295 1.980 4.785 2.100 ;
        RECT  4.665 0.960 4.735 1.080 ;
        RECT  4.545 0.960 4.665 1.790 ;
        RECT  4.425 0.650 4.590 0.770 ;
        RECT  4.305 0.650 4.425 1.860 ;
        RECT  4.295 0.380 4.415 0.530 ;
        RECT  3.720 0.650 4.305 0.770 ;
        RECT  2.770 1.740 4.305 1.860 ;
        RECT  3.690 0.410 4.295 0.530 ;
        RECT  3.740 1.070 4.185 1.330 ;
        RECT  3.620 0.890 3.740 1.620 ;
        RECT  3.570 0.380 3.690 0.530 ;
        RECT  3.600 0.890 3.620 1.010 ;
        RECT  3.130 1.500 3.620 1.620 ;
        RECT  3.480 0.650 3.600 1.010 ;
        RECT  3.295 0.380 3.570 0.500 ;
        RECT  3.250 1.190 3.500 1.310 ;
        RECT  3.420 0.650 3.480 0.770 ;
        RECT  2.900 0.620 3.420 0.770 ;
        RECT  3.035 0.350 3.295 0.500 ;
        RECT  3.035 1.980 3.295 2.190 ;
        RECT  3.120 1.060 3.250 1.310 ;
        RECT  2.475 1.060 3.120 1.180 ;
        RECT  2.710 0.380 3.035 0.500 ;
        RECT  2.205 1.980 3.035 2.100 ;
        RECT  2.650 1.340 2.770 1.860 ;
        RECT  2.590 0.380 2.710 0.540 ;
        RECT  1.655 0.420 2.590 0.540 ;
        RECT  2.375 0.660 2.475 1.570 ;
        RECT  2.355 0.660 2.375 1.810 ;
        RECT  1.805 0.660 2.355 0.780 ;
        RECT  2.255 1.450 2.355 1.810 ;
        RECT  2.045 1.690 2.255 1.810 ;
        RECT  2.075 1.980 2.205 2.140 ;
        RECT  1.845 2.020 2.075 2.140 ;
        RECT  1.775 1.380 1.895 1.900 ;
        RECT  1.650 2.020 1.845 2.190 ;
        RECT  1.655 1.380 1.775 1.500 ;
        RECT  1.535 0.420 1.655 1.500 ;
        RECT  1.530 1.725 1.650 2.190 ;
        RECT  0.645 1.725 1.530 1.845 ;
        RECT  0.975 1.425 1.000 1.595 ;
        RECT  0.855 0.680 0.975 1.595 ;
        RECT  0.830 1.020 0.855 1.595 ;
        RECT  0.715 1.020 0.830 1.280 ;
        RECT  0.595 0.705 0.645 0.875 ;
        RECT  0.595 1.445 0.645 2.135 ;
        RECT  0.475 0.705 0.595 2.135 ;
    END
END DFFNHX2AD
MACRO DFFNHX4AD
    CLASS CORE ;
    FOREIGN DFFNHX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.735 1.750 7.965 1.900 ;
        RECT  7.735 0.735 7.820 0.905 ;
        RECT  7.605 0.735 7.735 1.900 ;
        RECT  7.425 1.750 7.605 1.900 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.810 1.005 8.890 1.515 ;
        RECT  8.680 0.410 8.810 2.090 ;
        RECT  8.605 0.410 8.680 0.840 ;
        RECT  8.605 1.400 8.680 2.090 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.170 0.910 2.495 1.225 ;
        END
        AntennaGateArea 0.143 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.455 1.045 1.610 1.375 ;
        RECT  1.375 1.045 1.455 1.305 ;
        END
        AntennaGateArea 0.165 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.135 -0.210 9.240 0.210 ;
        RECT  8.965 -0.210 9.135 0.810 ;
        RECT  8.390 -0.210 8.965 0.210 ;
        RECT  8.270 -0.210 8.390 0.805 ;
        RECT  7.475 -0.210 8.270 0.210 ;
        RECT  7.215 -0.210 7.475 0.300 ;
        RECT  6.670 -0.210 7.215 0.210 ;
        RECT  6.410 -0.210 6.670 0.260 ;
        RECT  5.000 -0.210 6.410 0.210 ;
        RECT  4.740 -0.210 5.000 0.260 ;
        RECT  3.075 -0.210 4.740 0.210 ;
        RECT  2.555 -0.210 3.075 0.260 ;
        RECT  1.660 -0.210 2.555 0.210 ;
        RECT  1.490 -0.210 1.660 0.380 ;
        RECT  0.565 -0.210 1.490 0.210 ;
        RECT  0.395 -0.210 0.565 0.710 ;
        RECT  0.000 -0.210 0.395 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.135 2.310 9.240 2.730 ;
        RECT  8.965 1.680 9.135 2.730 ;
        RECT  8.345 2.310 8.965 2.730 ;
        RECT  8.175 2.265 8.345 2.730 ;
        RECT  7.540 2.310 8.175 2.730 ;
        RECT  7.370 2.265 7.540 2.730 ;
        RECT  6.790 2.310 7.370 2.730 ;
        RECT  6.530 2.220 6.790 2.730 ;
        RECT  5.150 2.310 6.530 2.730 ;
        RECT  4.980 2.265 5.150 2.730 ;
        RECT  4.205 2.310 4.980 2.730 ;
        RECT  3.945 2.290 4.205 2.730 ;
        RECT  3.015 2.310 3.945 2.730 ;
        RECT  2.755 2.260 3.015 2.730 ;
        RECT  1.615 2.310 2.755 2.730 ;
        RECT  1.355 2.010 1.615 2.730 ;
        RECT  0.615 2.310 1.355 2.730 ;
        RECT  0.445 1.750 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.240 2.520 ;
        LAYER M1 ;
        RECT  8.300 0.990 8.560 1.250 ;
        RECT  8.180 0.990 8.300 2.140 ;
        RECT  7.110 2.020 8.180 2.140 ;
        RECT  7.940 0.420 8.060 1.545 ;
        RECT  7.460 0.420 7.940 0.540 ;
        RECT  7.855 1.375 7.940 1.545 ;
        RECT  7.340 0.420 7.460 1.575 ;
        RECT  6.990 1.750 7.110 2.140 ;
        RECT  6.985 0.380 7.105 1.620 ;
        RECT  6.865 1.750 6.990 1.900 ;
        RECT  5.720 0.380 6.985 0.500 ;
        RECT  6.745 0.690 6.865 1.900 ;
        RECT  5.965 1.480 6.745 1.600 ;
        RECT  6.155 1.780 6.325 1.950 ;
        RECT  5.520 0.620 6.290 0.740 ;
        RECT  5.640 1.780 6.155 1.900 ;
        RECT  5.900 1.480 5.965 1.650 ;
        RECT  5.760 0.865 5.900 1.650 ;
        RECT  5.560 2.020 5.820 2.190 ;
        RECT  5.640 0.865 5.760 0.985 ;
        RECT  5.460 0.330 5.720 0.500 ;
        RECT  5.520 1.690 5.640 1.900 ;
        RECT  3.455 2.020 5.560 2.140 ;
        RECT  5.400 0.620 5.520 1.900 ;
        RECT  4.415 0.380 5.460 0.500 ;
        RECT  5.220 0.620 5.400 0.790 ;
        RECT  5.110 1.780 5.400 1.900 ;
        RECT  4.870 0.950 5.265 1.070 ;
        RECT  4.990 1.215 5.110 1.900 ;
        RECT  3.050 1.780 4.990 1.900 ;
        RECT  4.750 0.900 4.870 1.660 ;
        RECT  4.455 0.900 4.750 1.020 ;
        RECT  3.390 1.540 4.750 1.660 ;
        RECT  4.495 1.160 4.615 1.420 ;
        RECT  3.785 1.300 4.495 1.420 ;
        RECT  4.335 0.640 4.455 1.020 ;
        RECT  3.895 0.360 4.415 0.500 ;
        RECT  3.660 0.640 4.335 0.760 ;
        RECT  1.925 0.380 3.895 0.500 ;
        RECT  3.325 1.265 3.785 1.420 ;
        RECT  3.195 2.020 3.455 2.190 ;
        RECT  3.205 0.660 3.325 1.420 ;
        RECT  2.755 0.660 3.205 0.780 ;
        RECT  2.125 2.020 3.195 2.140 ;
        RECT  2.930 1.190 3.050 1.900 ;
        RECT  2.655 0.660 2.755 1.570 ;
        RECT  2.635 0.660 2.655 1.810 ;
        RECT  2.085 0.660 2.635 0.780 ;
        RECT  2.535 1.450 2.635 1.810 ;
        RECT  2.325 1.690 2.535 1.810 ;
        RECT  2.055 1.380 2.175 1.900 ;
        RECT  1.930 2.020 2.125 2.190 ;
        RECT  1.925 1.380 2.055 1.500 ;
        RECT  1.810 1.725 1.930 2.190 ;
        RECT  1.805 0.380 1.925 1.500 ;
        RECT  0.975 1.725 1.810 1.845 ;
        RECT  1.255 1.425 1.280 1.595 ;
        RECT  1.110 0.680 1.255 1.595 ;
        RECT  0.380 1.090 1.110 1.210 ;
        RECT  0.925 1.725 0.975 2.085 ;
        RECT  0.875 0.350 0.925 0.780 ;
        RECT  0.805 1.405 0.925 2.085 ;
        RECT  0.755 0.350 0.875 0.970 ;
        RECT  0.255 1.405 0.805 1.525 ;
        RECT  0.205 0.850 0.755 0.970 ;
        RECT  0.205 1.405 0.255 1.930 ;
        RECT  0.085 0.850 0.205 1.930 ;
    END
END DFFNHX4AD
MACRO DFFNHX8AD
    CLASS CORE ;
    FOREIGN DFFNHX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.720 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.595 0.660 11.690 0.830 ;
        RECT  11.595 1.780 11.680 1.900 ;
        RECT  11.465 0.660 11.595 1.900 ;
        RECT  11.420 1.330 11.465 1.900 ;
        RECT  11.085 1.330 11.420 1.780 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.275 1.000 13.510 1.625 ;
        RECT  13.105 0.380 13.275 2.145 ;
        RECT  13.025 0.665 13.105 1.625 ;
        RECT  12.555 0.665 13.025 0.915 ;
        RECT  12.555 1.375 13.025 1.625 ;
        RECT  12.385 0.410 12.555 0.915 ;
        RECT  12.385 1.375 12.555 2.155 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.570 1.125 3.885 1.295 ;
        RECT  3.150 1.125 3.570 1.375 ;
        END
        AntennaGateArea 0.262 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.080 2.090 1.250 ;
        RECT  1.750 1.080 1.890 1.655 ;
        END
        AntennaGateArea 0.275 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.635 -0.210 13.720 0.210 ;
        RECT  13.465 -0.210 13.635 0.810 ;
        RECT  12.915 -0.210 13.465 0.210 ;
        RECT  12.745 -0.210 12.915 0.490 ;
        RECT  12.170 -0.210 12.745 0.210 ;
        RECT  12.050 -0.210 12.170 0.805 ;
        RECT  11.355 -0.210 12.050 0.210 ;
        RECT  11.095 -0.210 11.355 0.260 ;
        RECT  8.420 -0.210 11.095 0.210 ;
        RECT  8.250 -0.210 8.420 0.260 ;
        RECT  7.660 -0.210 8.250 0.210 ;
        RECT  7.490 -0.210 7.660 0.260 ;
        RECT  6.860 -0.210 7.490 0.210 ;
        RECT  6.600 -0.210 6.860 0.260 ;
        RECT  4.795 -0.210 6.600 0.210 ;
        RECT  4.275 -0.210 4.795 0.260 ;
        RECT  3.550 -0.210 4.275 0.210 ;
        RECT  3.290 -0.210 3.550 0.380 ;
        RECT  1.995 -0.210 3.290 0.210 ;
        RECT  1.995 0.625 2.000 0.795 ;
        RECT  1.830 -0.210 1.995 0.795 ;
        RECT  1.825 -0.210 1.830 0.775 ;
        RECT  1.055 -0.210 1.825 0.210 ;
        RECT  0.885 -0.210 1.055 0.845 ;
        RECT  0.335 -0.210 0.885 0.210 ;
        RECT  0.165 -0.210 0.335 0.845 ;
        RECT  0.000 -0.210 0.165 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.635 2.310 13.720 2.730 ;
        RECT  13.465 1.775 13.635 2.730 ;
        RECT  12.915 2.310 13.465 2.730 ;
        RECT  12.745 1.765 12.915 2.730 ;
        RECT  12.125 2.310 12.745 2.730 ;
        RECT  11.955 2.265 12.125 2.730 ;
        RECT  11.255 2.310 11.955 2.730 ;
        RECT  11.085 2.265 11.255 2.730 ;
        RECT  8.145 2.310 11.085 2.730 ;
        RECT  7.885 2.005 8.145 2.730 ;
        RECT  7.405 2.310 7.885 2.730 ;
        RECT  7.145 2.265 7.405 2.730 ;
        RECT  5.860 2.310 7.145 2.730 ;
        RECT  5.600 2.290 5.860 2.730 ;
        RECT  4.420 2.310 5.600 2.730 ;
        RECT  4.160 2.260 4.420 2.730 ;
        RECT  3.550 2.310 4.160 2.730 ;
        RECT  3.290 2.020 3.550 2.730 ;
        RECT  2.065 2.310 3.290 2.730 ;
        RECT  1.805 2.190 2.065 2.730 ;
        RECT  1.000 2.310 1.805 2.730 ;
        RECT  0.830 1.630 1.000 2.730 ;
        RECT  0.280 2.310 0.830 2.730 ;
        RECT  0.110 1.630 0.280 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 13.720 2.520 ;
        LAYER M1 ;
        RECT  12.185 1.090 12.845 1.210 ;
        RECT  12.065 1.090 12.185 2.140 ;
        RECT  10.700 2.020 12.065 2.140 ;
        RECT  11.810 0.345 11.930 1.590 ;
        RECT  11.580 0.345 11.810 0.540 ;
        RECT  11.740 1.330 11.810 1.590 ;
        RECT  11.325 0.420 11.580 0.540 ;
        RECT  11.155 0.420 11.325 1.140 ;
        RECT  10.880 0.380 11.000 1.225 ;
        RECT  6.040 0.380 10.880 0.500 ;
        RECT  10.765 1.105 10.880 1.225 ;
        RECT  10.645 1.105 10.765 1.555 ;
        RECT  10.590 0.660 10.760 0.985 ;
        RECT  10.525 1.755 10.700 2.140 ;
        RECT  10.525 0.865 10.590 0.985 ;
        RECT  10.405 0.865 10.525 2.140 ;
        RECT  8.435 0.620 10.465 0.740 ;
        RECT  9.040 0.865 10.405 0.985 ;
        RECT  9.995 2.020 10.405 2.140 ;
        RECT  10.165 1.505 10.285 1.815 ;
        RECT  8.435 1.505 10.165 1.625 ;
        RECT  9.735 1.745 9.995 2.140 ;
        RECT  9.270 1.745 9.735 1.865 ;
        RECT  9.010 1.745 9.270 2.125 ;
        RECT  8.460 1.755 8.720 2.190 ;
        RECT  7.240 1.755 8.460 1.875 ;
        RECT  8.315 0.620 8.435 1.625 ;
        RECT  7.065 0.620 8.315 0.740 ;
        RECT  6.935 1.505 8.315 1.625 ;
        RECT  6.565 1.025 8.040 1.195 ;
        RECT  7.120 1.755 7.240 2.140 ;
        RECT  5.035 2.020 7.120 2.140 ;
        RECT  6.765 1.505 6.935 1.900 ;
        RECT  4.695 1.780 6.765 1.900 ;
        RECT  6.445 0.900 6.565 1.660 ;
        RECT  5.995 0.900 6.445 1.020 ;
        RECT  4.970 1.540 6.445 1.660 ;
        RECT  6.190 1.160 6.310 1.420 ;
        RECT  5.330 1.300 6.190 1.420 ;
        RECT  5.520 0.360 6.040 0.500 ;
        RECT  5.835 0.640 5.995 1.020 ;
        RECT  5.275 0.640 5.835 0.760 ;
        RECT  4.180 0.380 5.520 0.500 ;
        RECT  4.940 1.210 5.330 1.420 ;
        RECT  4.775 2.020 5.035 2.190 ;
        RECT  4.820 0.735 4.940 1.420 ;
        RECT  4.225 0.740 4.820 0.860 ;
        RECT  4.450 2.020 4.775 2.140 ;
        RECT  4.575 1.150 4.695 1.900 ;
        RECT  4.330 1.780 4.450 2.140 ;
        RECT  2.885 1.780 4.330 1.900 ;
        RECT  4.105 0.740 4.225 1.660 ;
        RECT  3.970 0.380 4.180 0.620 ;
        RECT  2.910 0.740 4.105 0.860 ;
        RECT  2.910 1.540 4.105 1.660 ;
        RECT  2.335 0.500 3.970 0.620 ;
        RECT  2.675 1.780 2.885 2.020 ;
        RECT  1.295 1.900 2.675 2.020 ;
        RECT  2.480 1.410 2.650 1.625 ;
        RECT  2.335 1.410 2.480 1.530 ;
        RECT  2.215 0.500 2.335 1.530 ;
        RECT  1.495 0.405 1.615 1.730 ;
        RECT  0.800 1.000 1.495 1.260 ;
        RECT  1.145 1.390 1.295 2.020 ;
        RECT  0.680 1.390 1.145 1.510 ;
        RECT  0.640 0.385 0.680 1.510 ;
        RECT  0.550 0.385 0.640 1.975 ;
        RECT  0.470 1.390 0.550 1.975 ;
    END
END DFFNHX8AD
MACRO DFFNSRHX1AD
    CLASS CORE ;
    FOREIGN DFFNSRHX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 1.080 3.025 1.375 ;
        END
        AntennaGateArea 0.115 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.225 1.020 7.345 1.280 ;
        RECT  5.855 1.080 7.225 1.200 ;
        RECT  5.625 1.080 5.855 1.330 ;
        END
        AntennaGateArea 0.108 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.510 1.425 8.635 1.710 ;
        RECT  8.390 0.910 8.510 1.710 ;
        RECT  8.170 0.910 8.390 1.030 ;
        END
        AntennaDiffArea 0.192 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.570 0.645 9.730 1.915 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.920 1.895 1.375 ;
        END
        AntennaGateArea 0.061 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.955 0.490 1.375 ;
        END
        AntennaGateArea 0.118 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.380 -0.210 9.800 0.210 ;
        RECT  9.120 -0.210 9.380 0.310 ;
        RECT  8.730 -0.210 9.120 0.210 ;
        RECT  8.470 -0.210 8.730 0.310 ;
        RECT  7.990 -0.210 8.470 0.210 ;
        RECT  7.730 -0.210 7.990 0.310 ;
        RECT  6.085 -0.210 7.730 0.210 ;
        RECT  5.825 -0.210 6.085 0.310 ;
        RECT  4.780 -0.210 5.825 0.210 ;
        RECT  4.520 -0.210 4.780 0.310 ;
        RECT  3.035 -0.210 4.520 0.210 ;
        RECT  2.775 -0.210 3.035 0.230 ;
        RECT  1.655 -0.210 2.775 0.210 ;
        RECT  1.535 -0.210 1.655 0.350 ;
        RECT  0.660 -0.210 1.535 0.210 ;
        RECT  0.490 -0.210 0.660 0.260 ;
        RECT  0.000 -0.210 0.490 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.315 2.310 9.800 2.730 ;
        RECT  8.885 2.150 9.315 2.730 ;
        RECT  7.530 2.310 8.885 2.730 ;
        RECT  7.270 2.230 7.530 2.730 ;
        RECT  5.915 2.310 7.270 2.730 ;
        RECT  5.655 2.290 5.915 2.730 ;
        RECT  5.285 2.310 5.655 2.730 ;
        RECT  5.025 2.220 5.285 2.730 ;
        RECT  4.345 2.310 5.025 2.730 ;
        RECT  4.085 2.220 4.345 2.730 ;
        RECT  2.840 2.310 4.085 2.730 ;
        RECT  2.320 2.220 2.840 2.730 ;
        RECT  1.840 2.310 2.320 2.730 ;
        RECT  1.670 2.220 1.840 2.730 ;
        RECT  0.560 2.310 1.670 2.730 ;
        RECT  0.390 1.925 0.560 2.730 ;
        RECT  0.000 2.310 0.390 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.800 2.520 ;
        LAYER M1 ;
        RECT  9.285 1.065 9.450 1.235 ;
        RECT  9.165 0.430 9.285 2.030 ;
        RECT  8.370 0.430 9.165 0.550 ;
        RECT  9.020 1.065 9.165 1.235 ;
        RECT  8.430 1.910 9.165 2.030 ;
        RECT  8.875 0.670 9.045 0.905 ;
        RECT  8.875 1.410 9.045 1.580 ;
        RECT  8.755 0.670 8.875 1.580 ;
        RECT  8.630 0.670 8.755 1.260 ;
        RECT  7.830 0.670 8.630 0.790 ;
        RECT  8.170 1.910 8.430 2.045 ;
        RECT  8.110 0.380 8.370 0.550 ;
        RECT  8.150 1.150 8.270 1.780 ;
        RECT  6.675 1.925 8.170 2.045 ;
        RECT  7.590 1.150 8.150 1.270 ;
        RECT  7.045 0.430 8.110 0.550 ;
        RECT  7.750 1.390 8.010 1.580 ;
        RECT  7.710 0.670 7.830 0.960 ;
        RECT  6.955 1.460 7.750 1.580 ;
        RECT  7.470 0.780 7.590 1.270 ;
        RECT  6.755 0.780 7.470 0.900 ;
        RECT  6.875 0.355 7.045 0.550 ;
        RECT  6.835 1.460 6.955 1.800 ;
        RECT  6.385 1.680 6.835 1.800 ;
        RECT  6.635 0.430 6.755 0.900 ;
        RECT  6.465 0.430 6.635 0.550 ;
        RECT  6.125 1.440 6.555 1.560 ;
        RECT  6.295 2.020 6.555 2.180 ;
        RECT  5.350 0.705 6.515 0.875 ;
        RECT  6.205 0.340 6.465 0.550 ;
        RECT  6.265 1.680 6.385 1.870 ;
        RECT  5.715 2.020 6.295 2.140 ;
        RECT  5.815 1.730 6.265 1.870 ;
        RECT  4.160 0.430 6.205 0.550 ;
        RECT  6.005 1.440 6.125 1.610 ;
        RECT  5.350 1.490 6.005 1.610 ;
        RECT  4.795 1.730 5.815 1.850 ;
        RECT  5.595 1.980 5.715 2.140 ;
        RECT  4.765 1.980 5.595 2.100 ;
        RECT  5.230 0.705 5.350 1.610 ;
        RECT  4.915 1.395 5.230 1.515 ;
        RECT  5.015 0.675 5.095 0.795 ;
        RECT  4.895 0.675 5.015 1.275 ;
        RECT  2.585 0.675 4.895 0.795 ;
        RECT  4.795 1.155 4.895 1.275 ;
        RECT  4.675 1.155 4.795 1.850 ;
        RECT  4.505 1.980 4.765 2.185 ;
        RECT  4.555 0.915 4.745 1.035 ;
        RECT  4.435 0.915 4.555 1.850 ;
        RECT  3.405 1.980 4.505 2.100 ;
        RECT  3.715 0.915 4.435 1.035 ;
        RECT  3.645 1.550 4.435 1.670 ;
        RECT  3.900 0.330 4.160 0.550 ;
        RECT  2.645 0.430 3.900 0.550 ;
        RECT  3.525 1.550 3.645 1.810 ;
        RECT  3.405 1.000 3.435 1.260 ;
        RECT  3.285 1.000 3.405 2.100 ;
        RECT  1.435 1.980 3.285 2.100 ;
        RECT  2.135 1.740 3.165 1.860 ;
        RECT  2.525 0.380 2.645 0.550 ;
        RECT  2.465 0.675 2.585 1.620 ;
        RECT  1.895 0.380 2.525 0.500 ;
        RECT  2.320 1.500 2.465 1.620 ;
        RECT  2.135 0.640 2.315 0.760 ;
        RECT  2.015 0.640 2.135 1.860 ;
        RECT  1.775 0.380 1.895 0.740 ;
        RECT  1.025 0.620 1.775 0.740 ;
        RECT  1.435 0.860 1.505 0.980 ;
        RECT  1.315 0.860 1.435 2.100 ;
        RECT  1.245 0.860 1.315 1.385 ;
        RECT  0.785 0.380 1.275 0.500 ;
        RECT  1.155 1.125 1.245 1.385 ;
        RECT  1.025 1.770 1.165 2.030 ;
        RECT  0.905 0.620 1.025 2.030 ;
        RECT  0.665 0.380 0.785 0.835 ;
        RECT  0.270 0.715 0.665 0.835 ;
        RECT  0.220 0.665 0.270 0.835 ;
        RECT  0.220 1.495 0.270 1.665 ;
        RECT  0.100 0.665 0.220 1.665 ;
    END
END DFFNSRHX1AD
MACRO DFFNSRHX2AD
    CLASS CORE ;
    FOREIGN DFFNSRHX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.010 3.110 1.375 ;
        END
        AntennaGateArea 0.137 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.225 1.020 7.345 1.280 ;
        RECT  5.855 1.080 7.225 1.200 ;
        RECT  5.625 1.080 5.855 1.330 ;
        END
        AntennaGateArea 0.134 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.510 1.425 8.635 1.710 ;
        RECT  8.390 0.910 8.510 1.710 ;
        RECT  8.170 0.910 8.390 1.030 ;
        END
        AntennaDiffArea 0.192 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.570 0.330 9.730 1.915 ;
        END
        AntennaDiffArea 0.368 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.920 1.895 1.375 ;
        END
        AntennaGateArea 0.088 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.040 0.770 1.375 ;
        END
        AntennaGateArea 0.127 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.330 -0.210 9.800 0.210 ;
        RECT  9.070 -0.210 9.330 0.310 ;
        RECT  8.730 -0.210 9.070 0.210 ;
        RECT  8.470 -0.210 8.730 0.310 ;
        RECT  7.990 -0.210 8.470 0.210 ;
        RECT  7.730 -0.210 7.990 0.310 ;
        RECT  6.085 -0.210 7.730 0.210 ;
        RECT  5.825 -0.210 6.085 0.310 ;
        RECT  4.780 -0.210 5.825 0.210 ;
        RECT  4.520 -0.210 4.780 0.310 ;
        RECT  2.985 -0.210 4.520 0.210 ;
        RECT  2.465 -0.210 2.985 0.230 ;
        RECT  1.920 -0.210 2.465 0.210 ;
        RECT  1.660 -0.210 1.920 0.315 ;
        RECT  0.545 -0.210 1.660 0.210 ;
        RECT  0.425 -0.210 0.545 0.400 ;
        RECT  0.000 -0.210 0.425 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.295 2.310 9.800 2.730 ;
        RECT  8.865 2.165 9.295 2.730 ;
        RECT  7.530 2.310 8.865 2.730 ;
        RECT  7.270 2.290 7.530 2.730 ;
        RECT  5.915 2.310 7.270 2.730 ;
        RECT  5.655 2.290 5.915 2.730 ;
        RECT  5.195 2.310 5.655 2.730 ;
        RECT  4.935 2.290 5.195 2.730 ;
        RECT  4.345 2.310 4.935 2.730 ;
        RECT  4.085 2.220 4.345 2.730 ;
        RECT  2.840 2.310 4.085 2.730 ;
        RECT  2.320 2.220 2.840 2.730 ;
        RECT  1.935 2.310 2.320 2.730 ;
        RECT  1.675 2.240 1.935 2.730 ;
        RECT  0.560 2.310 1.675 2.730 ;
        RECT  0.390 1.975 0.560 2.730 ;
        RECT  0.000 2.310 0.390 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.800 2.520 ;
        LAYER M1 ;
        RECT  9.285 1.065 9.450 1.235 ;
        RECT  9.165 0.430 9.285 2.045 ;
        RECT  8.370 0.430 9.165 0.550 ;
        RECT  9.020 1.065 9.165 1.235 ;
        RECT  8.170 1.910 9.165 2.045 ;
        RECT  8.875 0.670 9.045 0.905 ;
        RECT  8.875 1.410 9.045 1.580 ;
        RECT  8.755 0.670 8.875 1.580 ;
        RECT  8.630 0.670 8.755 1.260 ;
        RECT  7.830 0.670 8.630 0.790 ;
        RECT  8.110 0.380 8.370 0.550 ;
        RECT  8.150 1.150 8.270 1.780 ;
        RECT  6.675 1.925 8.170 2.045 ;
        RECT  7.590 1.150 8.150 1.270 ;
        RECT  7.045 0.430 8.110 0.550 ;
        RECT  7.750 1.390 8.010 1.580 ;
        RECT  7.710 0.670 7.830 0.960 ;
        RECT  6.955 1.460 7.750 1.580 ;
        RECT  7.470 0.780 7.590 1.270 ;
        RECT  6.755 0.780 7.470 0.900 ;
        RECT  6.875 0.355 7.045 0.550 ;
        RECT  6.835 1.460 6.955 1.800 ;
        RECT  6.385 1.680 6.835 1.800 ;
        RECT  6.635 0.435 6.755 0.900 ;
        RECT  6.465 0.435 6.635 0.555 ;
        RECT  6.125 1.440 6.555 1.560 ;
        RECT  5.350 0.705 6.515 0.875 ;
        RECT  6.205 0.330 6.465 0.555 ;
        RECT  6.265 1.680 6.385 1.880 ;
        RECT  6.095 2.020 6.355 2.190 ;
        RECT  5.825 1.730 6.265 1.880 ;
        RECT  4.160 0.435 6.205 0.555 ;
        RECT  6.005 1.440 6.125 1.610 ;
        RECT  5.715 2.020 6.095 2.140 ;
        RECT  5.350 1.490 6.005 1.610 ;
        RECT  4.795 1.730 5.825 1.850 ;
        RECT  5.595 1.980 5.715 2.140 ;
        RECT  4.765 1.980 5.595 2.100 ;
        RECT  5.230 0.705 5.350 1.610 ;
        RECT  4.915 1.395 5.230 1.515 ;
        RECT  5.015 0.675 5.095 0.795 ;
        RECT  4.895 0.675 5.015 1.275 ;
        RECT  2.600 0.675 4.895 0.795 ;
        RECT  4.795 1.155 4.895 1.275 ;
        RECT  4.675 1.155 4.795 1.850 ;
        RECT  4.505 1.980 4.765 2.185 ;
        RECT  4.555 0.915 4.745 1.035 ;
        RECT  4.435 0.915 4.555 1.850 ;
        RECT  3.405 1.980 4.505 2.100 ;
        RECT  3.715 0.915 4.435 1.035 ;
        RECT  3.645 1.550 4.435 1.670 ;
        RECT  3.900 0.330 4.160 0.555 ;
        RECT  1.895 0.435 3.900 0.555 ;
        RECT  3.525 1.550 3.645 1.810 ;
        RECT  3.405 1.000 3.435 1.260 ;
        RECT  3.285 1.000 3.405 2.100 ;
        RECT  1.435 1.980 3.285 2.100 ;
        RECT  2.135 1.740 3.165 1.860 ;
        RECT  2.480 0.675 2.600 1.620 ;
        RECT  2.320 1.500 2.480 1.620 ;
        RECT  2.135 0.765 2.330 0.885 ;
        RECT  2.015 0.765 2.135 1.860 ;
        RECT  1.775 0.435 1.895 0.740 ;
        RECT  1.025 0.620 1.775 0.740 ;
        RECT  0.785 0.380 1.540 0.500 ;
        RECT  1.435 0.860 1.505 0.980 ;
        RECT  1.315 0.860 1.435 2.100 ;
        RECT  1.245 0.860 1.315 1.385 ;
        RECT  1.145 1.125 1.245 1.385 ;
        RECT  1.025 1.760 1.165 2.020 ;
        RECT  0.905 0.620 1.025 2.020 ;
        RECT  0.665 0.380 0.785 0.835 ;
        RECT  0.270 0.715 0.665 0.835 ;
        RECT  0.220 0.665 0.270 0.835 ;
        RECT  0.220 1.510 0.270 1.680 ;
        RECT  0.100 0.665 0.220 1.680 ;
    END
END DFFNSRHX2AD
MACRO DFFNSRHX4AD
    CLASS CORE ;
    FOREIGN DFFNSRHX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.080 1.110 3.305 1.375 ;
        END
        AntennaGateArea 0.194 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.760 0.960 9.880 1.220 ;
        RECT  8.235 1.100 9.760 1.220 ;
        RECT  7.725 1.100 8.235 1.330 ;
        RECT  7.125 1.100 7.725 1.220 ;
        RECT  7.005 0.910 7.125 1.220 ;
        END
        AntennaGateArea 0.226 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.155 1.730 11.295 1.850 ;
        RECT  11.035 0.910 11.155 1.850 ;
        RECT  10.990 0.910 11.035 1.515 ;
        RECT  10.710 0.910 10.990 1.030 ;
        END
        AntennaDiffArea 0.198 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.435 1.005 12.530 1.515 ;
        RECT  12.265 0.365 12.435 2.175 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.920 2.275 1.375 ;
        END
        AntennaGateArea 0.153 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.110 0.770 1.375 ;
        END
        AntennaGateArea 0.167 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.795 -0.210 12.880 0.210 ;
        RECT  12.625 -0.210 12.795 0.795 ;
        RECT  12.050 -0.210 12.625 0.210 ;
        RECT  11.790 -0.210 12.050 0.310 ;
        RECT  11.370 -0.210 11.790 0.210 ;
        RECT  11.110 -0.210 11.370 0.310 ;
        RECT  10.500 -0.210 11.110 0.210 ;
        RECT  10.240 -0.210 10.500 0.310 ;
        RECT  8.250 -0.210 10.240 0.210 ;
        RECT  8.080 -0.210 8.250 0.260 ;
        RECT  6.980 -0.210 8.080 0.210 ;
        RECT  6.810 -0.210 6.980 0.260 ;
        RECT  6.125 -0.210 6.810 0.210 ;
        RECT  5.955 -0.210 6.125 0.255 ;
        RECT  5.235 -0.210 5.955 0.210 ;
        RECT  5.065 -0.210 5.235 0.255 ;
        RECT  3.275 -0.210 5.065 0.210 ;
        RECT  3.105 -0.210 3.275 0.255 ;
        RECT  1.895 -0.210 3.105 0.210 ;
        RECT  1.725 -0.210 1.895 0.450 ;
        RECT  0.610 -0.210 1.725 0.210 ;
        RECT  0.470 -0.210 0.610 0.750 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.795 2.310 12.880 2.730 ;
        RECT  12.625 1.635 12.795 2.730 ;
        RECT  12.075 2.310 12.625 2.730 ;
        RECT  11.905 1.960 12.075 2.730 ;
        RECT  11.695 2.310 11.905 2.730 ;
        RECT  11.435 2.210 11.695 2.730 ;
        RECT  10.020 2.310 11.435 2.730 ;
        RECT  9.760 2.220 10.020 2.730 ;
        RECT  7.380 2.310 9.760 2.730 ;
        RECT  7.210 2.260 7.380 2.730 ;
        RECT  6.450 2.310 7.210 2.730 ;
        RECT  6.280 2.260 6.450 2.730 ;
        RECT  4.995 2.310 6.280 2.730 ;
        RECT  4.825 2.260 4.995 2.730 ;
        RECT  3.340 2.310 4.825 2.730 ;
        RECT  2.820 2.260 3.340 2.730 ;
        RECT  2.280 2.310 2.820 2.730 ;
        RECT  2.020 2.290 2.280 2.730 ;
        RECT  1.520 2.310 2.020 2.730 ;
        RECT  1.260 2.290 1.520 2.730 ;
        RECT  0.575 2.310 1.260 2.730 ;
        RECT  0.405 2.105 0.575 2.730 ;
        RECT  0.000 2.310 0.405 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 12.880 2.520 ;
        LAYER M1 ;
        RECT  11.945 1.015 12.120 1.275 ;
        RECT  11.825 0.430 11.945 1.840 ;
        RECT  10.840 0.430 11.825 0.550 ;
        RECT  11.740 1.015 11.825 1.275 ;
        RECT  11.540 1.720 11.825 1.840 ;
        RECT  11.585 1.420 11.695 1.590 ;
        RECT  11.585 0.670 11.675 0.905 ;
        RECT  11.465 0.670 11.585 1.590 ;
        RECT  11.420 1.720 11.540 2.090 ;
        RECT  10.365 0.670 11.465 0.790 ;
        RECT  11.275 1.125 11.465 1.295 ;
        RECT  10.895 1.970 11.420 2.090 ;
        RECT  10.725 1.795 10.895 2.090 ;
        RECT  10.730 1.490 10.870 1.610 ;
        RECT  10.670 0.355 10.840 0.550 ;
        RECT  10.610 1.190 10.730 1.610 ;
        RECT  9.610 1.970 10.725 2.090 ;
        RECT  9.795 0.430 10.670 0.550 ;
        RECT  10.125 1.190 10.610 1.310 ;
        RECT  9.370 1.430 10.490 1.550 ;
        RECT  10.245 0.670 10.365 0.975 ;
        RECT  10.005 0.670 10.125 1.310 ;
        RECT  9.575 0.670 10.005 0.790 ;
        RECT  9.675 0.380 9.795 0.550 ;
        RECT  8.490 0.380 9.675 0.500 ;
        RECT  9.520 1.970 9.610 2.115 ;
        RECT  9.455 0.620 9.575 0.790 ;
        RECT  8.395 1.995 9.520 2.115 ;
        RECT  8.100 0.620 9.455 0.740 ;
        RECT  9.245 1.430 9.370 1.875 ;
        RECT  6.020 1.755 9.245 1.875 ;
        RECT  7.665 0.860 9.140 0.980 ;
        RECT  6.695 1.515 9.035 1.635 ;
        RECT  7.980 0.380 8.100 0.740 ;
        RECT  7.825 2.020 8.085 2.190 ;
        RECT  2.135 0.380 7.980 0.500 ;
        RECT  5.925 2.020 7.825 2.140 ;
        RECT  7.545 0.620 7.665 0.980 ;
        RECT  7.405 0.620 7.545 0.790 ;
        RECT  6.695 0.670 7.405 0.790 ;
        RECT  6.575 0.670 6.695 1.635 ;
        RECT  6.140 1.410 6.575 1.530 ;
        RECT  6.335 0.635 6.455 1.285 ;
        RECT  2.870 0.635 6.335 0.755 ;
        RECT  6.020 1.165 6.335 1.285 ;
        RECT  5.780 0.925 6.165 1.045 ;
        RECT  5.900 1.165 6.020 1.875 ;
        RECT  5.665 2.020 5.925 2.190 ;
        RECT  5.660 0.925 5.780 1.870 ;
        RECT  3.865 2.020 5.665 2.140 ;
        RECT  5.100 0.925 5.660 1.045 ;
        RECT  4.115 1.750 5.660 1.870 ;
        RECT  5.395 1.340 5.515 1.600 ;
        RECT  4.495 1.480 5.395 1.600 ;
        RECT  4.970 0.905 5.100 1.045 ;
        RECT  4.330 0.905 4.970 1.025 ;
        RECT  3.865 1.160 4.830 1.280 ;
        RECT  4.235 1.410 4.495 1.600 ;
        RECT  4.070 0.880 4.330 1.025 ;
        RECT  3.750 1.160 3.865 2.140 ;
        RECT  3.745 1.070 3.750 2.140 ;
        RECT  3.630 1.070 3.745 1.330 ;
        RECT  1.830 2.020 3.745 2.140 ;
        RECT  2.590 1.780 3.600 1.900 ;
        RECT  2.860 1.540 3.000 1.660 ;
        RECT  2.860 0.635 2.870 0.920 ;
        RECT  2.740 0.635 2.860 1.660 ;
        RECT  2.515 1.640 2.590 1.900 ;
        RECT  2.395 0.670 2.515 1.900 ;
        RECT  2.255 0.670 2.395 0.790 ;
        RECT  2.015 0.380 2.135 0.690 ;
        RECT  1.090 0.570 2.015 0.690 ;
        RECT  1.710 1.135 1.830 2.140 ;
        RECT  1.520 1.135 1.710 1.255 ;
        RECT  1.400 0.815 1.520 1.255 ;
        RECT  1.260 0.815 1.400 0.935 ;
        RECT  1.350 1.135 1.400 1.255 ;
        RECT  1.230 1.135 1.350 1.395 ;
        RECT  0.850 0.330 1.250 0.450 ;
        RECT  1.090 1.575 1.205 2.005 ;
        RECT  0.970 0.570 1.090 2.005 ;
        RECT  0.730 0.330 0.850 0.990 ;
        RECT  0.265 0.870 0.730 0.990 ;
        RECT  0.215 0.635 0.265 0.990 ;
        RECT  0.215 1.565 0.265 1.735 ;
        RECT  0.095 0.635 0.215 1.735 ;
    END
END DFFNSRHX4AD
MACRO DFFNSRHX8AD
    CLASS CORE ;
    FOREIGN DFFNSRHX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.350 1.070 3.585 1.375 ;
        END
        AntennaGateArea 0.235 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.995 0.925 10.115 1.220 ;
        RECT  8.515 1.100 9.995 1.220 ;
        RECT  8.005 1.100 8.515 1.330 ;
        RECT  7.390 1.100 8.005 1.220 ;
        RECT  7.220 0.965 7.390 1.220 ;
        END
        AntennaGateArea 0.262 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.550 1.730 11.685 1.850 ;
        RECT  11.425 0.910 11.550 1.850 ;
        RECT  11.130 0.910 11.425 1.515 ;
        RECT  11.095 0.910 11.130 1.030 ;
        END
        AntennaDiffArea 0.207 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.310 0.365 13.480 2.165 ;
        RECT  12.795 1.050 13.310 1.470 ;
        RECT  12.625 0.365 12.795 2.165 ;
        RECT  12.590 0.365 12.625 0.795 ;
        RECT  12.590 1.475 12.625 2.165 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.980 2.325 1.375 ;
        END
        AntennaGateArea 0.266 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.025 0.550 1.405 ;
        END
        AntennaGateArea 0.259 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.840 -0.210 14.000 0.210 ;
        RECT  13.670 -0.210 13.840 0.795 ;
        RECT  13.120 -0.210 13.670 0.210 ;
        RECT  12.950 -0.210 13.120 0.795 ;
        RECT  12.165 -0.210 12.950 0.210 ;
        RECT  11.645 -0.210 12.165 0.230 ;
        RECT  10.715 -0.210 11.645 0.210 ;
        RECT  10.455 -0.210 10.715 0.310 ;
        RECT  8.465 -0.210 10.455 0.210 ;
        RECT  8.345 -0.210 8.465 0.500 ;
        RECT  7.295 -0.210 8.345 0.210 ;
        RECT  7.035 -0.210 7.295 0.260 ;
        RECT  6.545 -0.210 7.035 0.210 ;
        RECT  6.025 -0.210 6.545 0.260 ;
        RECT  3.530 -0.210 6.025 0.210 ;
        RECT  3.270 -0.210 3.530 0.310 ;
        RECT  2.890 -0.210 3.270 0.210 ;
        RECT  2.630 -0.210 2.890 0.310 ;
        RECT  1.990 -0.210 2.630 0.210 ;
        RECT  1.730 -0.210 1.990 0.310 ;
        RECT  0.740 -0.210 1.730 0.210 ;
        RECT  0.480 -0.210 0.740 0.250 ;
        RECT  0.000 -0.210 0.480 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.840 2.310 14.000 2.730 ;
        RECT  13.670 1.475 13.840 2.730 ;
        RECT  13.120 2.310 13.670 2.730 ;
        RECT  12.950 1.735 13.120 2.730 ;
        RECT  12.375 2.310 12.950 2.730 ;
        RECT  11.855 2.220 12.375 2.730 ;
        RECT  10.330 2.310 11.855 2.730 ;
        RECT  10.070 2.220 10.330 2.730 ;
        RECT  7.775 2.310 10.070 2.730 ;
        RECT  7.515 2.260 7.775 2.730 ;
        RECT  6.845 2.310 7.515 2.730 ;
        RECT  6.585 2.260 6.845 2.730 ;
        RECT  5.375 2.310 6.585 2.730 ;
        RECT  5.115 2.260 5.375 2.730 ;
        RECT  3.410 2.310 5.115 2.730 ;
        RECT  2.890 2.260 3.410 2.730 ;
        RECT  1.475 2.310 2.890 2.730 ;
        RECT  1.305 2.185 1.475 2.730 ;
        RECT  0.565 2.310 1.305 2.730 ;
        RECT  0.395 2.265 0.565 2.730 ;
        RECT  0.000 2.310 0.395 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 14.000 2.520 ;
        LAYER M1 ;
        RECT  12.385 1.060 12.505 1.230 ;
        RECT  12.235 0.430 12.385 2.100 ;
        RECT  10.075 0.430 12.235 0.550 ;
        RECT  12.075 1.060 12.235 1.230 ;
        RECT  11.250 1.970 12.235 2.100 ;
        RECT  11.940 1.450 12.090 1.620 ;
        RECT  11.940 0.670 12.010 0.950 ;
        RECT  11.820 0.670 11.940 1.620 ;
        RECT  10.595 0.670 11.820 0.790 ;
        RECT  11.735 1.080 11.820 1.340 ;
        RECT  10.990 1.780 11.250 2.100 ;
        RECT  10.890 1.130 11.010 1.660 ;
        RECT  8.680 1.980 10.990 2.100 ;
        RECT  10.355 1.130 10.890 1.250 ;
        RECT  10.570 1.400 10.690 1.660 ;
        RECT  10.475 0.670 10.595 0.980 ;
        RECT  9.565 1.400 10.570 1.520 ;
        RECT  10.235 0.670 10.355 1.250 ;
        RECT  9.865 0.670 10.235 0.790 ;
        RECT  9.970 0.380 10.075 0.550 ;
        RECT  8.725 0.380 9.970 0.500 ;
        RECT  9.735 0.620 9.865 0.790 ;
        RECT  8.165 0.620 9.735 0.740 ;
        RECT  9.445 1.400 9.565 1.860 ;
        RECT  8.210 1.740 9.445 1.860 ;
        RECT  7.925 0.860 9.375 0.980 ;
        RECT  7.565 1.500 9.320 1.620 ;
        RECT  8.105 2.015 8.365 2.190 ;
        RECT  8.090 1.740 8.210 1.895 ;
        RECT  8.045 0.380 8.165 0.740 ;
        RECT  6.245 2.015 8.105 2.140 ;
        RECT  6.330 1.775 8.090 1.895 ;
        RECT  5.860 0.380 8.045 0.500 ;
        RECT  7.805 0.620 7.925 0.980 ;
        RECT  6.965 0.620 7.805 0.740 ;
        RECT  7.445 1.500 7.565 1.655 ;
        RECT  6.965 1.535 7.445 1.655 ;
        RECT  6.845 0.620 6.965 1.655 ;
        RECT  6.450 1.410 6.845 1.530 ;
        RECT  6.585 0.620 6.705 1.285 ;
        RECT  4.005 0.620 6.585 0.740 ;
        RECT  6.330 1.165 6.585 1.285 ;
        RECT  6.090 0.925 6.445 1.045 ;
        RECT  6.210 1.165 6.330 1.895 ;
        RECT  5.985 2.015 6.245 2.190 ;
        RECT  5.970 0.925 6.090 1.850 ;
        RECT  4.145 2.015 5.985 2.140 ;
        RECT  5.380 0.925 5.970 1.045 ;
        RECT  4.405 1.730 5.970 1.850 ;
        RECT  5.600 0.335 5.860 0.500 ;
        RECT  5.685 1.325 5.805 1.585 ;
        RECT  4.545 1.410 5.685 1.530 ;
        RECT  3.760 0.380 5.600 0.500 ;
        RECT  5.260 0.870 5.380 1.045 ;
        RECT  4.285 0.870 5.260 0.990 ;
        RECT  4.145 1.110 5.055 1.230 ;
        RECT  4.135 1.110 4.145 2.140 ;
        RECT  4.025 1.090 4.135 2.140 ;
        RECT  3.775 1.090 4.025 1.230 ;
        RECT  2.215 2.020 4.025 2.140 ;
        RECT  3.870 0.620 4.005 0.795 ;
        RECT  2.565 1.780 3.880 1.900 ;
        RECT  3.230 0.675 3.870 0.795 ;
        RECT  3.640 0.380 3.760 0.550 ;
        RECT  1.895 0.430 3.640 0.550 ;
        RECT  3.230 1.540 3.265 1.660 ;
        RECT  3.110 0.675 3.230 1.660 ;
        RECT  2.960 0.675 3.110 0.935 ;
        RECT  3.005 1.540 3.110 1.660 ;
        RECT  2.445 0.670 2.565 1.900 ;
        RECT  2.250 0.670 2.445 0.790 ;
        RECT  2.095 1.925 2.215 2.140 ;
        RECT  1.830 1.925 2.095 2.045 ;
        RECT  1.775 0.430 1.895 0.740 ;
        RECT  1.710 1.225 1.830 2.045 ;
        RECT  1.050 0.620 1.775 0.740 ;
        RECT  1.490 1.225 1.710 1.345 ;
        RECT  1.230 0.860 1.490 1.345 ;
        RECT  0.245 0.380 1.310 0.500 ;
        RECT  0.980 1.225 1.230 1.345 ;
        RECT  1.035 1.575 1.205 2.005 ;
        RECT  0.930 0.620 1.050 0.950 ;
        RECT  0.790 1.575 1.035 1.695 ;
        RECT  0.790 0.830 0.930 0.950 ;
        RECT  0.670 0.830 0.790 1.695 ;
        RECT  0.215 1.515 0.265 1.945 ;
        RECT  0.215 0.380 0.245 0.900 ;
        RECT  0.095 0.380 0.215 1.945 ;
    END
END DFFNSRHX8AD
MACRO DFFQX1AD
    CLASS CORE ;
    FOREIGN DFFQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.515 0.555 5.530 1.600 ;
        RECT  5.390 0.555 5.515 1.885 ;
        RECT  5.345 0.555 5.390 0.725 ;
        RECT  5.345 1.455 5.390 1.885 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.900 0.210 1.550 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.375 1.375 1.710 1.495 ;
        RECT  1.145 1.375 1.375 1.610 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.155 -0.210 5.600 0.210 ;
        RECT  5.155 0.560 5.200 0.680 ;
        RECT  4.985 -0.210 5.155 0.680 ;
        RECT  4.435 -0.210 4.985 0.210 ;
        RECT  4.940 0.560 4.985 0.680 ;
        RECT  4.265 -0.210 4.435 0.815 ;
        RECT  3.210 -0.210 4.265 0.210 ;
        RECT  3.040 -0.210 3.210 0.735 ;
        RECT  2.055 -0.210 3.040 0.210 ;
        RECT  1.885 -0.210 2.055 0.460 ;
        RECT  1.425 -0.210 1.885 0.210 ;
        RECT  1.255 -0.210 1.425 0.515 ;
        RECT  0.390 -0.210 1.255 0.210 ;
        RECT  0.130 -0.210 0.390 0.300 ;
        RECT  0.000 -0.210 0.130 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.155 2.310 5.600 2.730 ;
        RECT  4.985 1.520 5.155 2.730 ;
        RECT  4.415 2.310 4.985 2.730 ;
        RECT  4.245 1.550 4.415 2.730 ;
        RECT  3.210 2.310 4.245 2.730 ;
        RECT  2.950 2.160 3.210 2.730 ;
        RECT  2.150 2.310 2.950 2.730 ;
        RECT  1.890 2.160 2.150 2.730 ;
        RECT  1.385 2.310 1.890 2.730 ;
        RECT  1.215 2.105 1.385 2.730 ;
        RECT  0.285 2.310 1.215 2.730 ;
        RECT  0.115 2.085 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  5.080 0.800 5.200 1.400 ;
        RECT  4.800 0.800 5.080 0.920 ;
        RECT  4.775 1.280 5.080 1.400 ;
        RECT  3.825 1.040 4.960 1.160 ;
        RECT  4.630 0.645 4.800 0.920 ;
        RECT  4.605 1.280 4.775 1.745 ;
        RECT  4.080 1.280 4.605 1.400 ;
        RECT  3.760 0.350 4.020 0.500 ;
        RECT  3.655 0.645 3.825 1.800 ;
        RECT  3.535 0.380 3.760 0.500 ;
        RECT  3.535 1.920 3.730 2.165 ;
        RECT  3.470 0.380 3.535 2.165 ;
        RECT  3.415 0.380 3.470 2.040 ;
        RECT  2.965 0.890 3.415 1.010 ;
        RECT  1.710 1.920 3.415 2.040 ;
        RECT  3.175 1.130 3.295 1.785 ;
        RECT  2.440 1.665 3.175 1.785 ;
        RECT  2.800 0.890 2.965 1.250 ;
        RECT  2.680 0.590 2.885 0.710 ;
        RECT  2.680 1.415 2.825 1.535 ;
        RECT  2.560 0.330 2.680 1.535 ;
        RECT  2.420 0.330 2.560 0.450 ;
        RECT  2.320 0.690 2.440 1.785 ;
        RECT  1.955 1.665 2.320 1.785 ;
        RECT  2.080 0.895 2.200 1.370 ;
        RECT  0.795 0.895 2.080 1.015 ;
        RECT  1.835 1.135 1.955 1.785 ;
        RECT  1.050 0.655 1.850 0.775 ;
        RECT  1.040 1.135 1.835 1.255 ;
        RECT  1.570 1.635 1.710 2.155 ;
        RECT  0.990 1.865 1.570 1.985 ;
        RECT  0.930 0.420 1.050 0.775 ;
        RECT  0.730 1.865 0.990 2.110 ;
        RECT  0.480 0.420 0.930 0.540 ;
        RECT  0.745 0.675 0.795 1.015 ;
        RECT  0.745 1.575 0.795 1.745 ;
        RECT  0.625 0.675 0.745 1.745 ;
        RECT  0.480 1.865 0.730 1.985 ;
        RECT  0.360 0.420 0.480 1.985 ;
    END
END DFFQX1AD
MACRO DFFQX2AD
    CLASS CORE ;
    FOREIGN DFFQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.515 1.140 5.530 1.375 ;
        RECT  5.345 0.395 5.515 2.000 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.945 0.280 1.375 ;
        RECT  0.070 1.145 0.115 1.375 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.425 1.365 1.820 1.610 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.155 -0.210 5.600 0.210 ;
        RECT  4.985 -0.210 5.155 0.465 ;
        RECT  4.595 -0.210 4.985 0.210 ;
        RECT  4.425 -0.210 4.595 0.370 ;
        RECT  3.265 -0.210 4.425 0.210 ;
        RECT  3.005 -0.210 3.265 0.725 ;
        RECT  2.090 -0.210 3.005 0.210 ;
        RECT  1.920 -0.210 2.090 0.460 ;
        RECT  1.450 -0.210 1.920 0.210 ;
        RECT  1.280 -0.210 1.450 0.515 ;
        RECT  0.260 -0.210 1.280 0.210 ;
        RECT  0.090 -0.210 0.260 0.415 ;
        RECT  0.000 -0.210 0.090 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.155 2.310 5.600 2.730 ;
        RECT  4.985 1.975 5.155 2.730 ;
        RECT  4.570 2.310 4.985 2.730 ;
        RECT  4.310 1.510 4.570 2.730 ;
        RECT  3.265 2.310 4.310 2.730 ;
        RECT  3.005 2.190 3.265 2.730 ;
        RECT  2.185 2.310 3.005 2.730 ;
        RECT  1.925 2.190 2.185 2.730 ;
        RECT  1.410 2.310 1.925 2.730 ;
        RECT  1.240 2.145 1.410 2.730 ;
        RECT  0.260 2.310 1.240 2.730 ;
        RECT  0.090 2.105 0.260 2.730 ;
        RECT  0.000 2.310 0.090 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  4.930 0.630 5.050 1.390 ;
        RECT  4.715 0.630 4.930 0.800 ;
        RECT  4.885 1.270 4.930 1.390 ;
        RECT  4.715 1.270 4.885 1.625 ;
        RECT  4.570 1.030 4.810 1.150 ;
        RECT  4.330 1.270 4.715 1.390 ;
        RECT  4.450 0.625 4.570 1.150 ;
        RECT  3.850 0.625 4.450 0.745 ;
        RECT  4.210 1.020 4.330 1.390 ;
        RECT  3.610 1.950 4.100 2.070 ;
        RECT  3.815 0.330 4.075 0.500 ;
        RECT  3.730 0.625 3.850 1.620 ;
        RECT  3.505 0.380 3.815 0.500 ;
        RECT  3.625 0.625 3.730 0.745 ;
        RECT  3.505 0.865 3.610 2.070 ;
        RECT  3.490 0.380 3.505 2.070 ;
        RECT  3.385 0.380 3.490 0.985 ;
        RECT  1.805 1.950 3.490 2.070 ;
        RECT  2.965 0.865 3.385 0.985 ;
        RECT  3.310 1.105 3.360 1.275 ;
        RECT  3.190 1.105 3.310 1.830 ;
        RECT  2.480 1.710 3.190 1.830 ;
        RECT  2.845 0.865 2.965 1.255 ;
        RECT  2.720 1.430 2.885 1.550 ;
        RECT  2.720 0.565 2.830 0.735 ;
        RECT  2.600 0.330 2.720 1.550 ;
        RECT  2.395 0.330 2.600 0.450 ;
        RECT  2.360 0.570 2.480 1.830 ;
        RECT  2.310 0.570 2.360 0.740 ;
        RECT  1.095 1.125 2.360 1.245 ;
        RECT  2.265 1.710 2.360 1.830 ;
        RECT  0.820 0.885 2.220 1.005 ;
        RECT  1.080 0.645 1.875 0.765 ;
        RECT  1.545 1.745 1.805 2.125 ;
        RECT  1.015 1.875 1.545 1.995 ;
        RECT  0.960 0.410 1.080 0.765 ;
        RECT  0.755 1.875 1.015 2.115 ;
        RECT  0.520 0.410 0.960 0.530 ;
        RECT  0.700 0.675 0.820 1.755 ;
        RECT  0.520 1.875 0.755 1.995 ;
        RECT  0.650 0.675 0.700 0.845 ;
        RECT  0.650 1.585 0.700 1.755 ;
        RECT  0.400 0.410 0.520 1.995 ;
    END
END DFFQX2AD
MACRO DFFQX4AD
    CLASS CORE ;
    FOREIGN DFFQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.555 1.005 6.730 1.515 ;
        RECT  6.385 0.390 6.555 2.065 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.225 0.945 0.345 1.465 ;
        RECT  0.070 1.145 0.225 1.375 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.705 1.140 1.990 1.395 ;
        END
        AntennaGateArea 0.091 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.915 -0.210 7.000 0.210 ;
        RECT  6.745 -0.210 6.915 0.820 ;
        RECT  6.165 -0.210 6.745 0.210 ;
        RECT  5.995 -0.210 6.165 0.415 ;
        RECT  5.595 -0.210 5.995 0.210 ;
        RECT  5.425 -0.210 5.595 0.390 ;
        RECT  4.695 -0.210 5.425 0.210 ;
        RECT  4.525 -0.210 4.695 0.440 ;
        RECT  3.460 -0.210 4.525 0.210 ;
        RECT  3.200 -0.210 3.460 0.300 ;
        RECT  2.510 -0.210 3.200 0.210 ;
        RECT  2.250 -0.210 2.510 0.300 ;
        RECT  1.790 -0.210 2.250 0.210 ;
        RECT  1.530 -0.210 1.790 0.300 ;
        RECT  0.265 -0.210 1.530 0.210 ;
        RECT  0.095 -0.210 0.265 0.645 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.915 2.310 7.000 2.730 ;
        RECT  6.745 1.660 6.915 2.730 ;
        RECT  6.195 2.310 6.745 2.730 ;
        RECT  6.025 1.695 6.195 2.730 ;
        RECT  5.455 2.310 6.025 2.730 ;
        RECT  5.285 2.040 5.455 2.730 ;
        RECT  4.495 2.310 5.285 2.730 ;
        RECT  4.325 1.860 4.495 2.730 ;
        RECT  3.290 2.310 4.325 2.730 ;
        RECT  3.030 2.230 3.290 2.730 ;
        RECT  2.230 2.310 3.030 2.730 ;
        RECT  1.970 2.230 2.230 2.730 ;
        RECT  1.500 2.310 1.970 2.730 ;
        RECT  1.240 2.230 1.500 2.730 ;
        RECT  0.265 2.310 1.240 2.730 ;
        RECT  0.095 1.725 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.140 0.635 6.260 1.520 ;
        RECT  5.755 0.635 6.140 0.805 ;
        RECT  5.845 1.400 6.140 1.520 ;
        RECT  5.340 1.045 5.985 1.215 ;
        RECT  5.675 1.400 5.845 1.915 ;
        RECT  5.165 1.795 5.675 1.915 ;
        RECT  5.200 0.650 5.340 1.670 ;
        RECT  4.040 0.650 5.200 0.790 ;
        RECT  3.885 1.530 5.200 1.670 ;
        RECT  4.995 1.795 5.165 2.160 ;
        RECT  4.960 0.910 5.080 1.400 ;
        RECT  4.905 2.040 4.995 2.160 ;
        RECT  3.530 1.280 4.960 1.400 ;
        RECT  3.770 0.980 4.830 1.100 ;
        RECT  3.900 0.530 4.040 0.790 ;
        RECT  3.715 1.530 3.885 2.000 ;
        RECT  3.650 0.420 3.770 1.100 ;
        RECT  3.050 0.420 3.650 0.540 ;
        RECT  3.410 0.800 3.530 2.110 ;
        RECT  3.210 0.800 3.410 0.920 ;
        RECT  1.795 1.990 3.410 2.110 ;
        RECT  3.170 1.040 3.290 1.870 ;
        RECT  3.090 0.660 3.210 0.920 ;
        RECT  2.475 1.750 3.170 1.870 ;
        RECT  2.970 0.330 3.050 0.540 ;
        RECT  2.850 0.330 2.970 1.630 ;
        RECT  2.790 0.330 2.850 0.540 ;
        RECT  2.640 1.510 2.850 1.630 ;
        RECT  2.420 0.420 2.790 0.540 ;
        RECT  2.610 0.660 2.730 1.380 ;
        RECT  2.475 1.260 2.610 1.380 ;
        RECT  2.305 1.260 2.475 1.870 ;
        RECT  2.300 0.420 2.420 0.780 ;
        RECT  2.140 0.900 2.400 1.140 ;
        RECT  1.550 1.515 2.305 1.635 ;
        RECT  1.230 0.660 2.300 0.780 ;
        RECT  0.585 0.420 2.170 0.540 ;
        RECT  1.480 0.900 2.140 1.020 ;
        RECT  1.625 1.760 1.795 2.110 ;
        RECT  1.040 1.990 1.625 2.110 ;
        RECT  1.290 1.390 1.550 1.635 ;
        RECT  1.360 0.900 1.480 1.240 ;
        RECT  0.970 1.120 1.360 1.240 ;
        RECT  1.110 0.660 1.230 1.000 ;
        RECT  0.780 1.990 1.040 2.190 ;
        RECT  0.850 0.660 0.970 1.850 ;
        RECT  0.705 1.680 0.850 1.850 ;
        RECT  0.585 1.990 0.780 2.110 ;
        RECT  0.585 0.840 0.700 1.100 ;
        RECT  0.465 0.420 0.585 2.110 ;
    END
END DFFQX4AD
MACRO DFFQXLAD
    CLASS CORE ;
    FOREIGN DFFQXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.110 0.375 5.250 2.050 ;
        RECT  5.055 0.375 5.110 0.545 ;
        RECT  5.055 1.880 5.110 2.050 ;
        END
        AntennaDiffArea 0.138 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.900 0.210 1.550 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.375 1.375 1.715 1.495 ;
        RECT  1.145 1.375 1.375 1.610 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.865 -0.210 5.320 0.210 ;
        RECT  4.695 -0.210 4.865 0.545 ;
        RECT  4.435 -0.210 4.695 0.210 ;
        RECT  4.265 -0.210 4.435 0.815 ;
        RECT  3.255 -0.210 4.265 0.210 ;
        RECT  2.995 -0.210 3.255 0.770 ;
        RECT  2.055 -0.210 2.995 0.210 ;
        RECT  1.885 -0.210 2.055 0.460 ;
        RECT  1.425 -0.210 1.885 0.210 ;
        RECT  1.255 -0.210 1.425 0.515 ;
        RECT  0.255 -0.210 1.255 0.210 ;
        RECT  0.085 -0.210 0.255 0.360 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.865 2.310 5.320 2.730 ;
        RECT  4.695 1.890 4.865 2.730 ;
        RECT  4.415 2.310 4.695 2.730 ;
        RECT  4.245 1.550 4.415 2.730 ;
        RECT  3.210 2.310 4.245 2.730 ;
        RECT  2.950 2.190 3.210 2.730 ;
        RECT  2.150 2.310 2.950 2.730 ;
        RECT  1.890 2.190 2.150 2.730 ;
        RECT  1.375 2.310 1.890 2.730 ;
        RECT  1.205 2.115 1.375 2.730 ;
        RECT  0.285 2.310 1.205 2.730 ;
        RECT  0.115 2.085 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.320 2.520 ;
        LAYER M1 ;
        RECT  4.870 0.765 4.990 1.380 ;
        RECT  4.835 0.765 4.870 0.885 ;
        RECT  4.835 1.260 4.870 1.380 ;
        RECT  4.665 0.715 4.835 0.885 ;
        RECT  4.665 1.260 4.835 1.585 ;
        RECT  3.825 1.020 4.750 1.140 ;
        RECT  4.050 1.260 4.665 1.380 ;
        RECT  3.535 0.380 3.990 0.500 ;
        RECT  3.655 0.645 3.825 1.765 ;
        RECT  3.535 1.950 3.730 2.105 ;
        RECT  3.470 0.380 3.535 2.105 ;
        RECT  3.415 0.380 3.470 2.070 ;
        RECT  2.965 0.915 3.415 1.035 ;
        RECT  1.710 1.950 3.415 2.070 ;
        RECT  3.175 1.160 3.295 1.830 ;
        RECT  2.440 1.710 3.175 1.830 ;
        RECT  2.800 0.915 2.965 1.250 ;
        RECT  2.680 0.625 2.840 0.795 ;
        RECT  2.680 1.470 2.825 1.590 ;
        RECT  2.560 0.330 2.680 1.590 ;
        RECT  2.420 0.330 2.560 0.450 ;
        RECT  2.320 0.690 2.440 1.830 ;
        RECT  1.955 1.710 2.320 1.830 ;
        RECT  2.080 0.895 2.200 1.370 ;
        RECT  0.795 0.895 2.080 1.015 ;
        RECT  1.835 1.135 1.955 1.830 ;
        RECT  1.050 0.655 1.850 0.775 ;
        RECT  1.040 1.135 1.835 1.255 ;
        RECT  1.570 1.635 1.710 2.155 ;
        RECT  0.960 1.865 1.570 1.985 ;
        RECT  0.930 0.420 1.050 0.775 ;
        RECT  0.700 1.865 0.960 2.080 ;
        RECT  0.480 0.420 0.930 0.540 ;
        RECT  0.745 0.675 0.795 1.015 ;
        RECT  0.745 1.575 0.795 1.745 ;
        RECT  0.625 0.675 0.745 1.745 ;
        RECT  0.480 1.865 0.700 1.985 ;
        RECT  0.360 0.420 0.480 1.985 ;
    END
END DFFQXLAD
MACRO DFFRHQX1AD
    CLASS CORE ;
    FOREIGN DFFRHQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.640 1.460 5.780 1.580 ;
        RECT  5.520 1.280 5.640 1.580 ;
        RECT  4.790 1.280 5.520 1.400 ;
        RECT  4.505 1.100 4.790 1.400 ;
        END
        AntennaGateArea 0.097 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.330 0.655 7.490 1.920 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.685 0.900 1.870 1.160 ;
        RECT  1.470 0.865 1.685 1.160 ;
        END
        AntennaGateArea 0.075 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.445 1.050 0.770 1.375 ;
        END
        AntennaGateArea 0.114 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.045 -0.210 7.560 0.210 ;
        RECT  6.265 -0.210 7.045 0.325 ;
        RECT  4.735 -0.210 6.265 0.210 ;
        RECT  4.475 -0.210 4.735 0.300 ;
        RECT  3.690 -0.210 4.475 0.210 ;
        RECT  3.430 -0.210 3.690 0.300 ;
        RECT  2.325 -0.210 3.430 0.210 ;
        RECT  2.065 -0.210 2.325 0.300 ;
        RECT  1.770 -0.210 2.065 0.210 ;
        RECT  1.510 -0.210 1.770 0.300 ;
        RECT  0.690 -0.210 1.510 0.210 ;
        RECT  0.430 -0.210 0.690 0.300 ;
        RECT  0.000 -0.210 0.430 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.120 2.310 7.560 2.730 ;
        RECT  6.860 2.220 7.120 2.730 ;
        RECT  5.935 2.310 6.860 2.730 ;
        RECT  5.675 2.220 5.935 2.730 ;
        RECT  4.840 2.310 5.675 2.730 ;
        RECT  4.580 2.220 4.840 2.730 ;
        RECT  4.080 2.310 4.580 2.730 ;
        RECT  3.820 2.220 4.080 2.730 ;
        RECT  3.250 2.310 3.820 2.730 ;
        RECT  2.990 2.220 3.250 2.730 ;
        RECT  1.895 2.310 2.990 2.730 ;
        RECT  1.635 2.175 1.895 2.730 ;
        RECT  0.555 2.310 1.635 2.730 ;
        RECT  0.385 1.885 0.555 2.730 ;
        RECT  0.000 2.310 0.385 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  6.960 0.495 7.080 2.080 ;
        RECT  6.270 0.495 6.960 0.615 ;
        RECT  5.575 1.960 6.960 2.080 ;
        RECT  6.620 0.735 6.670 0.905 ;
        RECT  6.620 1.375 6.670 1.545 ;
        RECT  6.500 0.735 6.620 1.545 ;
        RECT  6.020 1.680 6.515 1.800 ;
        RECT  6.260 1.120 6.500 1.240 ;
        RECT  6.150 0.495 6.270 0.730 ;
        RECT  6.140 0.980 6.260 1.240 ;
        RECT  5.385 0.610 6.150 0.730 ;
        RECT  5.900 1.040 6.020 1.800 ;
        RECT  5.145 1.040 5.900 1.160 ;
        RECT  5.455 1.740 5.575 2.080 ;
        RECT  5.280 1.740 5.455 1.860 ;
        RECT  5.265 0.610 5.385 0.870 ;
        RECT  5.160 2.070 5.300 2.190 ;
        RECT  5.040 1.965 5.160 2.190 ;
        RECT  5.025 0.330 5.145 1.160 ;
        RECT  4.965 1.530 5.135 1.700 ;
        RECT  3.660 1.965 5.040 2.085 ;
        RECT  4.865 0.330 5.025 0.540 ;
        RECT  4.415 1.580 4.965 1.700 ;
        RECT  4.785 0.660 4.905 0.920 ;
        RECT  1.510 0.420 4.865 0.540 ;
        RECT  4.380 0.660 4.785 0.780 ;
        RECT  4.380 1.580 4.415 1.845 ;
        RECT  4.240 0.660 4.380 1.845 ;
        RECT  3.810 0.660 4.240 0.780 ;
        RECT  3.740 1.310 4.240 1.430 ;
        RECT  3.075 0.980 4.100 1.100 ;
        RECT  3.400 1.965 3.660 2.190 ;
        RECT  3.075 1.710 3.540 1.830 ;
        RECT  2.350 1.965 3.400 2.085 ;
        RECT  2.955 0.815 3.075 1.830 ;
        RECT  2.950 0.815 2.955 0.935 ;
        RECT  2.590 1.710 2.955 1.830 ;
        RECT  2.830 0.675 2.950 0.935 ;
        RECT  2.635 1.150 2.735 1.410 ;
        RECT  2.515 0.660 2.635 1.410 ;
        RECT  2.470 1.570 2.590 1.830 ;
        RECT  2.110 0.660 2.515 0.780 ;
        RECT  2.350 0.965 2.395 1.225 ;
        RECT  2.230 0.965 2.350 2.085 ;
        RECT  1.230 1.840 2.230 1.960 ;
        RECT  1.990 0.660 2.110 1.660 ;
        RECT  1.805 0.660 1.990 0.780 ;
        RECT  1.390 0.420 1.510 0.710 ;
        RECT  1.300 1.425 1.455 1.595 ;
        RECT  1.300 0.590 1.390 0.710 ;
        RECT  1.180 0.590 1.300 1.595 ;
        RECT  1.010 1.775 1.230 1.960 ;
        RECT  1.040 0.340 1.180 0.460 ;
        RECT  1.150 0.590 1.180 0.850 ;
        RECT  1.155 1.110 1.180 1.370 ;
        RECT  0.920 0.340 1.040 0.540 ;
        RECT  0.890 0.740 1.010 1.960 ;
        RECT  0.240 0.420 0.920 0.540 ;
        RECT  0.720 0.740 0.890 0.860 ;
        RECT  0.120 0.420 0.240 1.660 ;
    END
END DFFRHQX1AD
MACRO DFFRHQX2AD
    CLASS CORE ;
    FOREIGN DFFRHQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.800 1.175 5.920 1.635 ;
        RECT  5.050 1.175 5.800 1.295 ;
        RECT  4.830 1.000 5.050 1.375 ;
        END
        AntennaGateArea 0.141 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.330 0.385 7.490 2.020 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.005 1.955 1.265 ;
        RECT  1.725 1.005 1.890 1.760 ;
        END
        AntennaGateArea 0.077 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.050 0.530 1.655 ;
        END
        AntennaGateArea 0.119 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.090 -0.210 7.560 0.210 ;
        RECT  6.830 -0.210 7.090 0.310 ;
        RECT  6.520 -0.210 6.830 0.210 ;
        RECT  6.260 -0.210 6.520 0.310 ;
        RECT  4.790 -0.210 6.260 0.210 ;
        RECT  4.530 -0.210 4.790 0.260 ;
        RECT  3.800 -0.210 4.530 0.210 ;
        RECT  3.540 -0.210 3.800 0.260 ;
        RECT  2.455 -0.210 3.540 0.210 ;
        RECT  2.195 -0.210 2.455 0.260 ;
        RECT  1.860 -0.210 2.195 0.210 ;
        RECT  1.600 -0.210 1.860 0.260 ;
        RECT  0.680 -0.210 1.600 0.210 ;
        RECT  0.420 -0.210 0.680 0.310 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.140 2.310 7.560 2.730 ;
        RECT  6.880 1.995 7.140 2.730 ;
        RECT  6.170 2.310 6.880 2.730 ;
        RECT  6.140 2.210 6.170 2.730 ;
        RECT  5.875 2.185 6.140 2.730 ;
        RECT  4.870 2.310 5.875 2.730 ;
        RECT  4.700 2.265 4.870 2.730 ;
        RECT  4.240 2.310 4.700 2.730 ;
        RECT  3.980 2.220 4.240 2.730 ;
        RECT  3.420 2.310 3.980 2.730 ;
        RECT  3.160 2.220 3.420 2.730 ;
        RECT  1.880 2.310 3.160 2.730 ;
        RECT  1.620 2.220 1.880 2.730 ;
        RECT  0.520 2.310 1.620 2.730 ;
        RECT  0.380 1.900 0.520 2.730 ;
        RECT  0.000 2.310 0.380 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  6.970 0.520 7.090 1.875 ;
        RECT  5.530 0.520 6.970 0.640 ;
        RECT  5.520 1.755 6.970 1.875 ;
        RECT  6.780 0.760 6.850 0.880 ;
        RECT  6.660 0.760 6.780 1.590 ;
        RECT  6.590 0.760 6.660 1.140 ;
        RECT  6.400 1.020 6.590 1.140 ;
        RECT  6.390 1.370 6.510 1.630 ;
        RECT  6.280 0.950 6.400 1.210 ;
        RECT  6.160 1.370 6.390 1.490 ;
        RECT  6.040 0.935 6.160 1.490 ;
        RECT  5.290 0.935 6.040 1.055 ;
        RECT  5.410 0.520 5.530 0.780 ;
        RECT  5.280 1.440 5.420 1.560 ;
        RECT  5.170 0.380 5.290 1.055 ;
        RECT  5.160 1.440 5.280 1.720 ;
        RECT  3.340 0.380 5.170 0.500 ;
        RECT  4.640 1.600 5.160 1.720 ;
        RECT  5.040 1.930 5.160 2.190 ;
        RECT  4.870 0.650 5.040 0.820 ;
        RECT  3.790 1.970 5.040 2.090 ;
        RECT  4.640 0.700 4.870 0.820 ;
        RECT  4.595 0.700 4.640 1.820 ;
        RECT  4.520 0.700 4.595 1.845 ;
        RECT  3.915 0.700 4.520 0.820 ;
        RECT  4.425 1.600 4.520 1.845 ;
        RECT  3.260 1.260 4.400 1.380 ;
        RECT  3.795 0.700 3.915 1.140 ;
        RECT  3.420 1.020 3.795 1.140 ;
        RECT  3.530 1.910 3.790 2.090 ;
        RECT  3.260 1.560 3.670 1.680 ;
        RECT  2.460 1.970 3.530 2.090 ;
        RECT  3.080 0.345 3.340 0.500 ;
        RECT  3.135 0.715 3.260 1.680 ;
        RECT  2.900 0.715 3.135 0.835 ;
        RECT  2.720 1.560 3.135 1.680 ;
        RECT  1.410 0.380 3.080 0.500 ;
        RECT  2.770 0.955 2.870 1.215 ;
        RECT  2.650 0.660 2.770 1.215 ;
        RECT  2.600 1.400 2.720 1.680 ;
        RECT  2.220 0.660 2.650 0.780 ;
        RECT  2.460 0.995 2.490 1.255 ;
        RECT  2.340 0.995 2.460 2.090 ;
        RECT  1.230 1.970 2.340 2.090 ;
        RECT  2.100 0.660 2.220 1.745 ;
        RECT  1.915 0.660 2.100 0.865 ;
        RECT  1.410 1.465 1.455 1.635 ;
        RECT  1.275 0.380 1.410 1.635 ;
        RECT  0.890 1.135 1.275 1.395 ;
        RECT  0.970 1.850 1.230 2.090 ;
        RECT  0.895 0.410 1.155 0.615 ;
        RECT  0.770 1.850 0.970 1.970 ;
        RECT  0.770 0.735 0.935 0.905 ;
        RECT  0.230 0.495 0.895 0.615 ;
        RECT  0.650 0.735 0.770 1.970 ;
        RECT  0.110 0.495 0.230 1.715 ;
    END
END DFFRHQX2AD
MACRO DFFRHQX4AD
    CLASS CORE ;
    FOREIGN DFFRHQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.885 1.330 7.330 1.450 ;
        RECT  6.765 1.220 6.885 1.450 ;
        RECT  5.855 1.220 6.765 1.360 ;
        RECT  5.625 1.100 5.855 1.360 ;
        END
        AntennaGateArea 0.242 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.795 1.005 8.890 1.515 ;
        RECT  8.625 0.405 8.795 2.170 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.710 0.860 1.890 1.375 ;
        END
        AntennaGateArea 0.12 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.490 1.375 ;
        END
        AntennaGateArea 0.193 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.155 -0.210 9.240 0.210 ;
        RECT  8.985 -0.210 9.155 0.835 ;
        RECT  8.365 -0.210 8.985 0.210 ;
        RECT  8.195 -0.210 8.365 0.350 ;
        RECT  7.755 -0.210 8.195 0.210 ;
        RECT  7.585 -0.210 7.755 0.350 ;
        RECT  5.765 -0.210 7.585 0.210 ;
        RECT  5.595 -0.210 5.765 0.495 ;
        RECT  4.345 -0.210 5.595 0.210 ;
        RECT  4.085 -0.210 4.345 0.300 ;
        RECT  3.140 -0.210 4.085 0.210 ;
        RECT  2.880 -0.210 3.140 0.300 ;
        RECT  1.860 -0.210 2.880 0.210 ;
        RECT  1.600 -0.210 1.860 0.240 ;
        RECT  0.645 -0.210 1.600 0.210 ;
        RECT  0.475 -0.210 0.645 0.315 ;
        RECT  0.000 -0.210 0.475 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.155 2.310 9.240 2.730 ;
        RECT  8.985 1.730 9.155 2.730 ;
        RECT  8.425 2.310 8.985 2.730 ;
        RECT  8.255 2.020 8.425 2.730 ;
        RECT  7.425 2.310 8.255 2.730 ;
        RECT  7.255 2.010 7.425 2.730 ;
        RECT  5.635 2.310 7.255 2.730 ;
        RECT  5.465 2.250 5.635 2.730 ;
        RECT  4.870 2.310 5.465 2.730 ;
        RECT  4.610 2.250 4.870 2.730 ;
        RECT  3.630 2.310 4.610 2.730 ;
        RECT  3.370 2.250 3.630 2.730 ;
        RECT  2.210 2.310 3.370 2.730 ;
        RECT  1.950 1.990 2.210 2.730 ;
        RECT  1.490 2.310 1.950 2.730 ;
        RECT  1.230 1.990 1.490 2.730 ;
        RECT  0.565 2.310 1.230 2.730 ;
        RECT  0.395 2.030 0.565 2.730 ;
        RECT  0.000 2.310 0.395 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.240 2.520 ;
        LAYER M1 ;
        RECT  8.335 0.470 8.455 1.890 ;
        RECT  7.220 0.470 8.335 0.590 ;
        RECT  6.070 1.770 8.335 1.890 ;
        RECT  8.095 0.760 8.215 1.520 ;
        RECT  7.880 0.760 8.095 0.880 ;
        RECT  7.620 1.400 8.095 1.520 ;
        RECT  7.810 1.020 7.930 1.280 ;
        RECT  7.615 1.020 7.810 1.140 ;
        RECT  7.500 1.260 7.620 1.520 ;
        RECT  7.495 0.710 7.615 1.140 ;
        RECT  6.950 0.710 7.495 0.830 ;
        RECT  7.100 0.380 7.220 0.590 ;
        RECT  6.990 0.380 7.100 0.500 ;
        RECT  6.730 0.330 6.990 0.500 ;
        RECT  6.830 0.620 6.950 0.830 ;
        RECT  6.640 2.010 6.900 2.190 ;
        RECT  5.435 0.620 6.830 0.740 ;
        RECT  5.970 0.380 6.730 0.500 ;
        RECT  6.475 1.480 6.645 1.650 ;
        RECT  4.450 2.010 6.640 2.130 ;
        RECT  5.505 0.860 6.610 0.980 ;
        RECT  5.900 1.480 6.475 1.600 ;
        RECT  5.780 1.480 5.900 1.765 ;
        RECT  5.505 1.645 5.780 1.765 ;
        RECT  5.385 0.860 5.505 1.765 ;
        RECT  5.315 0.420 5.435 0.740 ;
        RECT  5.140 0.860 5.385 0.980 ;
        RECT  4.750 1.645 5.385 1.765 ;
        RECT  3.960 0.420 5.315 0.540 ;
        RECT  4.350 1.125 5.180 1.245 ;
        RECT  4.880 0.700 5.140 0.980 ;
        RECT  4.630 1.365 4.750 1.765 ;
        RECT  4.490 1.365 4.630 1.485 ;
        RECT  4.190 2.010 4.450 2.190 ;
        RECT  4.230 0.680 4.350 1.810 ;
        RECT  2.445 0.680 4.230 0.800 ;
        RECT  4.000 1.580 4.230 1.810 ;
        RECT  2.690 2.010 4.190 2.130 ;
        RECT  3.940 1.340 4.110 1.460 ;
        RECT  2.930 1.580 4.000 1.700 ;
        RECT  3.700 0.350 3.960 0.540 ;
        RECT  3.820 1.110 3.940 1.460 ;
        RECT  3.110 1.110 3.820 1.230 ;
        RECT  2.760 0.420 3.700 0.540 ;
        RECT  2.990 0.925 3.110 1.230 ;
        RECT  2.500 0.925 2.990 1.045 ;
        RECT  2.810 1.580 2.930 1.840 ;
        RECT  2.640 0.380 2.760 0.540 ;
        RECT  2.570 1.750 2.690 2.130 ;
        RECT  1.590 0.380 2.640 0.500 ;
        RECT  1.175 1.750 2.570 1.870 ;
        RECT  2.380 0.925 2.500 1.630 ;
        RECT  2.275 0.620 2.445 0.800 ;
        RECT  2.150 0.925 2.380 1.045 ;
        RECT  2.030 0.620 2.150 1.045 ;
        RECT  1.890 0.620 2.030 0.740 ;
        RECT  1.590 1.510 1.850 1.630 ;
        RECT  1.470 0.380 1.590 1.630 ;
        RECT  1.220 0.620 1.470 0.740 ;
        RECT  0.850 1.165 1.470 1.285 ;
        RECT  0.900 0.330 1.290 0.450 ;
        RECT  1.005 1.405 1.175 1.870 ;
        RECT  0.730 1.405 1.005 1.525 ;
        RECT  0.800 0.675 0.920 0.935 ;
        RECT  0.780 0.330 0.900 0.555 ;
        RECT  0.730 0.815 0.800 0.935 ;
        RECT  0.230 0.435 0.780 0.555 ;
        RECT  0.610 0.815 0.730 1.525 ;
        RECT  0.110 0.435 0.230 1.730 ;
    END
END DFFRHQX4AD
MACRO DFFRHQX8AD
    CLASS CORE ;
    FOREIGN DFFRHQX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.810 1.220 8.070 1.390 ;
        RECT  6.695 1.220 7.810 1.360 ;
        RECT  6.300 1.100 6.695 1.360 ;
        END
        AntennaGateArea 0.293 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.025 0.365 10.195 2.170 ;
        RECT  9.475 1.005 10.025 1.515 ;
        RECT  9.305 0.365 9.475 2.170 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.265 0.910 2.640 1.175 ;
        END
        AntennaGateArea 0.232 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.560 1.375 ;
        END
        AntennaGateArea 0.353 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.555 -0.210 10.640 0.210 ;
        RECT  10.385 -0.210 10.555 0.795 ;
        RECT  9.835 -0.210 10.385 0.210 ;
        RECT  9.665 -0.210 9.835 0.795 ;
        RECT  9.045 -0.210 9.665 0.210 ;
        RECT  8.875 -0.210 9.045 0.350 ;
        RECT  8.555 -0.210 8.875 0.210 ;
        RECT  8.385 -0.210 8.555 0.350 ;
        RECT  6.505 -0.210 8.385 0.210 ;
        RECT  6.335 -0.210 6.505 0.500 ;
        RECT  5.085 -0.210 6.335 0.210 ;
        RECT  4.825 -0.210 5.085 0.300 ;
        RECT  3.880 -0.210 4.825 0.210 ;
        RECT  3.620 -0.210 3.880 0.300 ;
        RECT  2.510 -0.210 3.620 0.210 ;
        RECT  2.250 -0.210 2.510 0.260 ;
        RECT  1.675 -0.210 2.250 0.210 ;
        RECT  1.675 0.330 1.725 0.500 ;
        RECT  1.555 -0.210 1.675 0.500 ;
        RECT  0.680 -0.210 1.555 0.210 ;
        RECT  0.420 -0.210 0.680 0.400 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.530 2.310 10.640 2.730 ;
        RECT  10.410 1.435 10.530 2.730 ;
        RECT  9.835 2.310 10.410 2.730 ;
        RECT  9.665 1.730 9.835 2.730 ;
        RECT  9.090 2.310 9.665 2.730 ;
        RECT  8.830 2.210 9.090 2.730 ;
        RECT  8.200 2.310 8.830 2.730 ;
        RECT  7.940 2.120 8.200 2.730 ;
        RECT  6.375 2.310 7.940 2.730 ;
        RECT  6.205 2.265 6.375 2.730 ;
        RECT  5.660 2.310 6.205 2.730 ;
        RECT  5.400 2.210 5.660 2.730 ;
        RECT  4.370 2.310 5.400 2.730 ;
        RECT  4.110 2.210 4.370 2.730 ;
        RECT  3.295 2.310 4.110 2.730 ;
        RECT  3.125 2.210 3.295 2.730 ;
        RECT  2.555 2.310 3.125 2.730 ;
        RECT  2.385 1.985 2.555 2.730 ;
        RECT  1.835 2.310 2.385 2.730 ;
        RECT  1.665 1.990 1.835 2.730 ;
        RECT  0.615 2.310 1.665 2.730 ;
        RECT  0.445 1.855 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.640 2.520 ;
        LAYER M1 ;
        RECT  9.065 0.470 9.185 2.000 ;
        RECT  8.025 0.470 9.065 0.590 ;
        RECT  7.935 1.880 9.065 2.000 ;
        RECT  8.790 0.760 8.910 1.520 ;
        RECT  8.590 0.760 8.790 0.880 ;
        RECT  8.430 1.400 8.790 1.520 ;
        RECT  8.550 1.020 8.670 1.280 ;
        RECT  8.355 1.020 8.550 1.140 ;
        RECT  8.310 1.400 8.430 1.760 ;
        RECT  8.235 0.710 8.355 1.140 ;
        RECT  8.190 1.500 8.310 1.760 ;
        RECT  7.690 0.710 8.235 0.830 ;
        RECT  7.905 0.380 8.025 0.590 ;
        RECT  7.815 1.770 7.935 2.000 ;
        RECT  7.710 0.380 7.905 0.500 ;
        RECT  6.770 1.770 7.815 1.890 ;
        RECT  7.450 0.330 7.710 0.500 ;
        RECT  7.570 0.620 7.690 0.830 ;
        RECT  7.380 2.010 7.640 2.190 ;
        RECT  6.175 0.620 7.570 0.740 ;
        RECT  6.885 0.380 7.450 0.500 ;
        RECT  7.215 1.480 7.385 1.650 ;
        RECT  6.665 2.010 7.380 2.130 ;
        RECT  6.160 0.860 7.325 0.980 ;
        RECT  6.640 1.480 7.215 1.600 ;
        RECT  6.715 0.330 6.885 0.500 ;
        RECT  6.545 1.970 6.665 2.130 ;
        RECT  6.520 1.480 6.640 1.765 ;
        RECT  5.190 1.970 6.545 2.090 ;
        RECT  6.160 1.645 6.520 1.765 ;
        RECT  6.055 0.420 6.175 0.740 ;
        RECT  6.040 0.860 6.160 1.765 ;
        RECT  4.700 0.420 6.055 0.540 ;
        RECT  5.880 0.860 6.040 0.980 ;
        RECT  5.490 1.645 6.040 1.765 ;
        RECT  5.090 1.125 5.920 1.245 ;
        RECT  5.620 0.700 5.880 0.980 ;
        RECT  5.370 1.365 5.490 1.765 ;
        RECT  5.230 1.365 5.370 1.485 ;
        RECT  4.930 1.970 5.190 2.190 ;
        RECT  4.970 0.680 5.090 1.845 ;
        RECT  4.400 0.680 4.970 0.800 ;
        RECT  3.670 1.725 4.970 1.845 ;
        RECT  3.305 1.970 4.930 2.090 ;
        RECT  4.690 1.320 4.850 1.440 ;
        RECT  4.440 0.350 4.700 0.540 ;
        RECT  4.560 1.110 4.690 1.440 ;
        RECT  3.850 1.110 4.560 1.230 ;
        RECT  3.455 0.420 4.440 0.540 ;
        RECT  4.280 0.670 4.400 0.800 ;
        RECT  3.185 0.670 4.280 0.790 ;
        RECT  3.730 0.920 3.850 1.230 ;
        RECT  2.915 0.920 3.730 1.040 ;
        RECT  3.550 1.585 3.670 1.845 ;
        RECT  3.305 1.255 3.610 1.375 ;
        RECT  3.335 0.380 3.455 0.540 ;
        RECT  2.440 0.380 3.335 0.500 ;
        RECT  3.185 1.255 3.305 2.090 ;
        RECT  3.015 0.620 3.185 0.790 ;
        RECT  1.200 1.745 3.185 1.865 ;
        RECT  2.880 0.920 2.915 1.625 ;
        RECT  2.795 0.620 2.880 1.625 ;
        RECT  2.760 0.620 2.795 1.040 ;
        RECT  2.745 1.455 2.795 1.625 ;
        RECT  2.675 0.620 2.760 0.790 ;
        RECT  2.320 0.380 2.440 0.740 ;
        RECT  2.145 0.620 2.320 0.740 ;
        RECT  2.145 1.455 2.195 1.625 ;
        RECT  2.025 0.620 2.145 1.625 ;
        RECT  1.320 0.620 2.025 0.740 ;
        RECT  1.175 0.330 1.435 0.500 ;
        RECT  1.200 0.620 1.320 1.400 ;
        RECT  1.010 1.280 1.200 1.400 ;
        RECT  1.080 1.620 1.200 2.140 ;
        RECT  0.920 0.380 1.175 0.500 ;
        RECT  0.890 1.620 1.080 1.740 ;
        RECT  0.890 0.760 1.060 0.880 ;
        RECT  0.800 0.380 0.920 0.640 ;
        RECT  0.770 0.760 0.890 1.740 ;
        RECT  0.230 0.520 0.800 0.640 ;
        RECT  0.110 0.330 0.230 1.965 ;
    END
END DFFRHQX8AD
MACRO DFFRQX1AD
    CLASS CORE ;
    FOREIGN DFFRQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.070 4.905 1.190 ;
        RECT  4.280 0.430 4.400 1.190 ;
        RECT  3.835 0.430 4.280 0.550 ;
        RECT  3.715 0.430 3.835 0.665 ;
        RECT  3.335 0.545 3.715 0.665 ;
        RECT  3.200 0.545 3.335 0.770 ;
        RECT  3.030 0.380 3.200 0.770 ;
        RECT  1.305 0.380 3.030 0.500 ;
        END
        AntennaGateArea 0.1 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.930 0.660 6.090 1.930 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.310 0.910 1.685 1.190 ;
        END
        AntennaGateArea 0.067 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.195 0.865 0.375 1.215 ;
        RECT  0.070 0.865 0.195 1.095 ;
        END
        AntennaGateArea 0.048 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 -0.210 6.160 0.210 ;
        RECT  5.545 -0.210 5.715 0.870 ;
        RECT  4.720 -0.210 5.545 0.210 ;
        RECT  4.550 -0.210 4.720 0.935 ;
        RECT  3.580 -0.210 4.550 0.210 ;
        RECT  3.320 -0.210 3.580 0.415 ;
        RECT  1.185 -0.210 3.320 0.210 ;
        RECT  1.025 -0.210 1.185 0.500 ;
        RECT  0.690 -0.210 1.025 0.210 ;
        RECT  0.430 -0.210 0.690 0.325 ;
        RECT  0.000 -0.210 0.430 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 2.310 6.160 2.730 ;
        RECT  5.545 1.410 5.715 2.730 ;
        RECT  4.850 2.310 5.545 2.730 ;
        RECT  4.680 1.855 4.850 2.730 ;
        RECT  3.130 2.310 4.680 2.730 ;
        RECT  2.960 1.830 3.130 2.730 ;
        RECT  1.510 2.310 2.960 2.730 ;
        RECT  1.250 2.015 1.510 2.730 ;
        RECT  0.700 2.310 1.250 2.730 ;
        RECT  0.440 1.685 0.700 2.730 ;
        RECT  0.000 2.310 0.440 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.415 1.000 5.810 1.260 ;
        RECT  5.295 0.755 5.415 1.735 ;
        RECT  5.135 0.755 5.295 0.875 ;
        RECT  4.525 1.615 5.295 1.735 ;
        RECT  5.055 0.995 5.175 1.455 ;
        RECT  4.060 1.335 5.055 1.455 ;
        RECT  4.355 1.615 4.525 2.165 ;
        RECT  3.940 1.925 4.200 2.110 ;
        RECT  4.060 0.765 4.110 0.935 ;
        RECT  3.940 0.765 4.060 1.755 ;
        RECT  3.780 1.635 3.940 1.755 ;
        RECT  3.370 1.925 3.940 2.045 ;
        RECT  3.610 0.790 3.795 0.910 ;
        RECT  3.490 0.790 3.610 1.805 ;
        RECT  2.970 1.185 3.490 1.305 ;
        RECT  3.250 1.580 3.370 2.045 ;
        RECT  2.705 1.580 3.250 1.700 ;
        RECT  2.850 1.185 2.970 1.445 ;
        RECT  2.585 0.620 2.705 1.700 ;
        RECT  2.505 1.930 2.625 2.190 ;
        RECT  1.940 0.620 2.585 0.740 ;
        RECT  2.495 1.170 2.585 1.430 ;
        RECT  2.330 1.930 2.505 2.050 ;
        RECT  2.330 0.875 2.465 1.045 ;
        RECT  2.210 0.875 2.330 2.050 ;
        RECT  1.120 1.775 2.210 1.895 ;
        RECT  1.820 0.620 1.940 1.445 ;
        RECT  1.090 1.325 1.820 1.445 ;
        RECT  0.860 1.775 1.120 1.955 ;
        RECT  0.995 1.325 1.090 1.530 ;
        RECT  0.875 0.620 0.995 1.530 ;
        RECT  0.765 0.620 0.875 0.790 ;
        RECT  0.830 1.410 0.875 1.530 ;
        RECT  0.625 0.995 0.730 1.255 ;
        RECT  0.505 0.625 0.625 1.565 ;
        RECT  0.265 0.625 0.505 0.745 ;
        RECT  0.265 1.445 0.505 1.565 ;
        RECT  0.095 0.575 0.265 0.745 ;
        RECT  0.095 1.445 0.265 1.615 ;
    END
END DFFRQX1AD
MACRO DFFRQX2AD
    CLASS CORE ;
    FOREIGN DFFRQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.070 4.905 1.190 ;
        RECT  4.280 0.430 4.400 1.190 ;
        RECT  3.835 0.430 4.280 0.550 ;
        RECT  3.715 0.430 3.835 0.665 ;
        RECT  3.335 0.545 3.715 0.665 ;
        RECT  3.200 0.545 3.335 0.770 ;
        RECT  3.030 0.380 3.200 0.770 ;
        RECT  1.305 0.380 3.030 0.500 ;
        END
        AntennaGateArea 0.106 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.930 0.335 6.090 1.930 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.310 0.910 1.685 1.190 ;
        END
        AntennaGateArea 0.067 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.195 0.865 0.375 1.215 ;
        RECT  0.070 0.865 0.195 1.095 ;
        END
        AntennaGateArea 0.048 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 -0.210 6.160 0.210 ;
        RECT  5.545 -0.210 5.715 0.810 ;
        RECT  4.720 -0.210 5.545 0.210 ;
        RECT  4.550 -0.210 4.720 0.935 ;
        RECT  3.580 -0.210 4.550 0.210 ;
        RECT  3.320 -0.210 3.580 0.415 ;
        RECT  1.185 -0.210 3.320 0.210 ;
        RECT  1.025 -0.210 1.185 0.500 ;
        RECT  0.690 -0.210 1.025 0.210 ;
        RECT  0.430 -0.210 0.690 0.325 ;
        RECT  0.000 -0.210 0.430 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 2.310 6.160 2.730 ;
        RECT  5.545 1.410 5.715 2.730 ;
        RECT  4.850 2.310 5.545 2.730 ;
        RECT  4.680 1.855 4.850 2.730 ;
        RECT  3.130 2.310 4.680 2.730 ;
        RECT  2.960 1.830 3.130 2.730 ;
        RECT  1.510 2.310 2.960 2.730 ;
        RECT  1.250 2.015 1.510 2.730 ;
        RECT  0.700 2.310 1.250 2.730 ;
        RECT  0.440 1.685 0.700 2.730 ;
        RECT  0.000 2.310 0.440 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.415 1.000 5.810 1.260 ;
        RECT  5.295 0.755 5.415 1.735 ;
        RECT  5.135 0.755 5.295 0.875 ;
        RECT  4.525 1.615 5.295 1.735 ;
        RECT  5.055 0.995 5.175 1.455 ;
        RECT  4.060 1.335 5.055 1.455 ;
        RECT  4.355 1.615 4.525 2.165 ;
        RECT  3.940 1.925 4.200 2.110 ;
        RECT  4.060 0.765 4.110 0.935 ;
        RECT  3.940 0.765 4.060 1.755 ;
        RECT  3.780 1.635 3.940 1.755 ;
        RECT  3.370 1.925 3.940 2.045 ;
        RECT  3.610 0.790 3.795 0.910 ;
        RECT  3.490 0.790 3.610 1.805 ;
        RECT  2.970 1.185 3.490 1.305 ;
        RECT  3.250 1.580 3.370 2.045 ;
        RECT  2.705 1.580 3.250 1.700 ;
        RECT  2.850 1.185 2.970 1.445 ;
        RECT  2.585 0.620 2.705 1.700 ;
        RECT  2.505 1.930 2.625 2.190 ;
        RECT  1.940 0.620 2.585 0.740 ;
        RECT  2.495 1.170 2.585 1.430 ;
        RECT  2.330 1.930 2.505 2.050 ;
        RECT  2.330 0.875 2.465 1.045 ;
        RECT  2.210 0.875 2.330 2.050 ;
        RECT  1.120 1.775 2.210 1.895 ;
        RECT  1.820 0.620 1.940 1.445 ;
        RECT  1.045 1.325 1.820 1.445 ;
        RECT  0.860 1.775 1.120 1.955 ;
        RECT  0.995 1.325 1.045 1.555 ;
        RECT  0.875 0.620 0.995 1.555 ;
        RECT  0.765 0.620 0.875 0.790 ;
        RECT  0.625 0.995 0.730 1.255 ;
        RECT  0.505 0.625 0.625 1.565 ;
        RECT  0.265 0.625 0.505 0.745 ;
        RECT  0.265 1.445 0.505 1.565 ;
        RECT  0.095 0.575 0.265 0.745 ;
        RECT  0.095 1.445 0.265 1.615 ;
    END
END DFFRQX2AD
MACRO DFFRQX4AD
    CLASS CORE ;
    FOREIGN DFFRQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.070 4.915 1.190 ;
        RECT  4.280 0.430 4.400 1.190 ;
        RECT  3.835 0.430 4.280 0.550 ;
        RECT  3.715 0.430 3.835 0.630 ;
        RECT  3.335 0.510 3.715 0.630 ;
        RECT  3.200 0.510 3.335 0.770 ;
        RECT  3.030 0.380 3.200 0.770 ;
        RECT  1.600 0.380 3.030 0.500 ;
        RECT  1.480 0.380 1.600 0.745 ;
        RECT  1.260 0.625 1.480 0.745 ;
        RECT  1.140 0.625 1.260 1.205 ;
        END
        AntennaGateArea 0.143 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.995 0.695 6.090 1.680 ;
        RECT  5.950 0.445 5.995 1.975 ;
        RECT  5.825 0.445 5.950 0.875 ;
        RECT  5.825 1.500 5.950 1.975 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 0.865 1.685 1.190 ;
        END
        AntennaGateArea 0.067 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.985 0.375 1.215 ;
        RECT  0.070 0.865 0.210 1.215 ;
        END
        AntennaGateArea 0.048 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.370 -0.210 6.440 0.210 ;
        RECT  6.210 -0.210 6.370 0.925 ;
        RECT  5.630 -0.210 6.210 0.210 ;
        RECT  5.460 -0.210 5.630 0.550 ;
        RECT  4.755 -0.210 5.460 0.210 ;
        RECT  4.555 -0.210 4.755 0.920 ;
        RECT  3.580 -0.210 4.555 0.210 ;
        RECT  3.320 -0.210 3.580 0.390 ;
        RECT  1.195 -0.210 3.320 0.210 ;
        RECT  1.025 -0.210 1.195 0.380 ;
        RECT  0.635 -0.210 1.025 0.210 ;
        RECT  0.465 -0.210 0.635 0.315 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.370 2.310 6.440 2.730 ;
        RECT  6.210 1.500 6.370 2.730 ;
        RECT  5.635 2.310 6.210 2.730 ;
        RECT  5.465 1.865 5.635 2.730 ;
        RECT  4.775 2.310 5.465 2.730 ;
        RECT  4.605 1.875 4.775 2.730 ;
        RECT  3.130 2.310 4.605 2.730 ;
        RECT  2.960 1.830 3.130 2.730 ;
        RECT  1.500 2.310 2.960 2.730 ;
        RECT  1.240 2.015 1.500 2.730 ;
        RECT  0.695 2.310 1.240 2.730 ;
        RECT  0.435 1.620 0.695 2.730 ;
        RECT  0.000 2.310 0.435 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.440 2.520 ;
        LAYER M1 ;
        RECT  5.560 1.000 5.820 1.260 ;
        RECT  5.440 0.725 5.560 1.735 ;
        RECT  5.180 0.725 5.440 0.895 ;
        RECT  4.460 1.615 5.440 1.735 ;
        RECT  5.140 1.185 5.260 1.455 ;
        RECT  4.110 1.335 5.140 1.455 ;
        RECT  4.340 1.615 4.460 2.190 ;
        RECT  3.930 1.925 4.190 2.110 ;
        RECT  3.940 0.735 4.110 1.780 ;
        RECT  3.825 1.610 3.940 1.780 ;
        RECT  3.370 1.925 3.930 2.045 ;
        RECT  3.610 0.760 3.795 0.880 ;
        RECT  3.490 0.760 3.610 1.805 ;
        RECT  2.825 1.270 3.490 1.390 ;
        RECT  3.250 1.535 3.370 2.045 ;
        RECT  2.705 1.535 3.250 1.655 ;
        RECT  2.585 0.620 2.705 1.655 ;
        RECT  2.505 1.775 2.625 2.190 ;
        RECT  1.940 0.620 2.585 0.740 ;
        RECT  2.495 1.170 2.585 1.430 ;
        RECT  2.375 1.775 2.505 1.895 ;
        RECT  2.375 0.875 2.465 1.045 ;
        RECT  2.255 0.875 2.375 1.895 ;
        RECT  1.120 1.775 2.255 1.895 ;
        RECT  1.820 0.620 1.940 1.445 ;
        RECT  1.045 1.325 1.820 1.445 ;
        RECT  0.860 1.775 1.120 1.955 ;
        RECT  0.995 1.325 1.045 1.555 ;
        RECT  0.875 0.575 0.995 1.555 ;
        RECT  0.765 0.575 0.875 0.745 ;
        RECT  0.625 0.995 0.730 1.255 ;
        RECT  0.505 0.625 0.625 1.495 ;
        RECT  0.255 0.625 0.505 0.745 ;
        RECT  0.255 1.375 0.505 1.495 ;
        RECT  0.085 0.575 0.255 0.745 ;
        RECT  0.085 1.375 0.255 1.545 ;
    END
END DFFRQX4AD
MACRO DFFRQXLAD
    CLASS CORE ;
    FOREIGN DFFRQXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.400 1.070 4.905 1.190 ;
        RECT  4.280 0.430 4.400 1.190 ;
        RECT  3.835 0.430 4.280 0.550 ;
        RECT  3.715 0.430 3.835 0.665 ;
        RECT  3.335 0.545 3.715 0.665 ;
        RECT  3.200 0.545 3.335 0.770 ;
        RECT  3.030 0.380 3.200 0.770 ;
        RECT  1.305 0.380 3.030 0.500 ;
        END
        AntennaGateArea 0.1 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.930 0.655 6.090 1.725 ;
        END
        AntennaDiffArea 0.138 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.310 0.910 1.685 1.190 ;
        END
        AntennaGateArea 0.067 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.195 0.865 0.375 1.215 ;
        RECT  0.070 0.865 0.195 1.095 ;
        END
        AntennaGateArea 0.048 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 -0.210 6.160 0.210 ;
        RECT  5.545 -0.210 5.715 0.870 ;
        RECT  4.720 -0.210 5.545 0.210 ;
        RECT  4.550 -0.210 4.720 0.935 ;
        RECT  3.580 -0.210 4.550 0.210 ;
        RECT  3.320 -0.210 3.580 0.415 ;
        RECT  1.185 -0.210 3.320 0.210 ;
        RECT  1.025 -0.210 1.185 0.500 ;
        RECT  0.690 -0.210 1.025 0.210 ;
        RECT  0.430 -0.210 0.690 0.325 ;
        RECT  0.000 -0.210 0.430 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 2.310 6.160 2.730 ;
        RECT  5.545 1.465 5.715 2.730 ;
        RECT  4.850 2.310 5.545 2.730 ;
        RECT  4.680 1.855 4.850 2.730 ;
        RECT  3.130 2.310 4.680 2.730 ;
        RECT  2.960 1.830 3.130 2.730 ;
        RECT  1.510 2.310 2.960 2.730 ;
        RECT  1.250 2.015 1.510 2.730 ;
        RECT  0.700 2.310 1.250 2.730 ;
        RECT  0.440 1.685 0.700 2.730 ;
        RECT  0.000 2.310 0.440 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.415 1.000 5.810 1.260 ;
        RECT  5.295 0.755 5.415 1.735 ;
        RECT  5.135 0.755 5.295 0.875 ;
        RECT  4.525 1.615 5.295 1.735 ;
        RECT  5.055 0.995 5.175 1.455 ;
        RECT  4.060 1.335 5.055 1.455 ;
        RECT  4.355 1.615 4.525 2.165 ;
        RECT  3.940 1.925 4.200 2.110 ;
        RECT  4.060 0.765 4.110 0.935 ;
        RECT  3.940 0.765 4.060 1.755 ;
        RECT  3.780 1.635 3.940 1.755 ;
        RECT  3.370 1.925 3.940 2.045 ;
        RECT  3.610 0.790 3.795 0.910 ;
        RECT  3.490 0.790 3.610 1.805 ;
        RECT  2.970 1.185 3.490 1.305 ;
        RECT  3.250 1.580 3.370 2.045 ;
        RECT  2.705 1.580 3.250 1.700 ;
        RECT  2.850 1.185 2.970 1.445 ;
        RECT  2.585 0.620 2.705 1.700 ;
        RECT  2.505 1.930 2.625 2.190 ;
        RECT  1.940 0.620 2.585 0.740 ;
        RECT  2.495 1.170 2.585 1.430 ;
        RECT  2.330 1.930 2.505 2.050 ;
        RECT  2.330 0.875 2.465 1.045 ;
        RECT  2.210 0.875 2.330 2.050 ;
        RECT  1.120 1.775 2.210 1.895 ;
        RECT  1.820 0.620 1.940 1.445 ;
        RECT  1.090 1.325 1.820 1.445 ;
        RECT  0.860 1.775 1.120 1.955 ;
        RECT  0.995 1.325 1.090 1.530 ;
        RECT  0.875 0.620 0.995 1.530 ;
        RECT  0.765 0.620 0.875 0.790 ;
        RECT  0.830 1.410 0.875 1.530 ;
        RECT  0.625 0.995 0.730 1.255 ;
        RECT  0.505 0.625 0.625 1.565 ;
        RECT  0.265 0.625 0.505 0.745 ;
        RECT  0.265 1.445 0.505 1.565 ;
        RECT  0.095 0.575 0.265 0.745 ;
        RECT  0.095 1.445 0.265 1.615 ;
    END
END DFFRQXLAD
MACRO DFFRX1AD
    CLASS CORE ;
    FOREIGN DFFRX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 0.400 5.160 1.140 ;
        RECT  3.815 0.400 5.040 0.520 ;
        RECT  3.695 0.400 3.815 0.760 ;
        RECT  3.590 0.640 3.695 0.760 ;
        RECT  3.470 0.640 3.590 1.220 ;
        RECT  3.335 0.640 3.470 0.760 ;
        RECT  3.215 0.380 3.335 0.760 ;
        RECT  2.020 0.380 3.215 0.500 ;
        RECT  1.900 0.380 2.020 0.540 ;
        RECT  1.050 0.420 1.900 0.540 ;
        RECT  0.870 0.420 1.050 0.880 ;
        END
        AntennaGateArea 0.102 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.940 0.585 6.090 0.865 ;
        RECT  5.820 0.585 5.940 1.590 ;
        END
        AntennaDiffArea 0.174 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.510 0.705 6.650 1.930 ;
        RECT  6.465 0.705 6.510 0.875 ;
        RECT  6.485 1.410 6.510 1.930 ;
        END
        AntennaDiffArea 0.203 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.240 0.230 1.655 ;
        END
        AntennaGateArea 0.067 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.910 1.655 1.060 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.290 -0.210 6.720 0.210 ;
        RECT  6.030 -0.210 6.290 0.355 ;
        RECT  5.060 -0.210 6.030 0.210 ;
        RECT  4.800 -0.210 5.060 0.280 ;
        RECT  3.575 -0.210 4.800 0.210 ;
        RECT  3.455 -0.210 3.575 0.475 ;
        RECT  1.780 -0.210 3.455 0.210 ;
        RECT  1.520 -0.210 1.780 0.300 ;
        RECT  1.240 -0.210 1.520 0.210 ;
        RECT  0.980 -0.210 1.240 0.300 ;
        RECT  0.000 -0.210 0.980 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.085 2.310 6.720 2.730 ;
        RECT  5.705 2.150 6.085 2.730 ;
        RECT  5.035 2.310 5.705 2.730 ;
        RECT  4.775 2.210 5.035 2.730 ;
        RECT  3.540 2.310 4.775 2.730 ;
        RECT  3.370 1.830 3.540 2.730 ;
        RECT  3.010 2.310 3.370 2.730 ;
        RECT  2.750 2.105 3.010 2.730 ;
        RECT  1.615 2.310 2.750 2.730 ;
        RECT  1.185 2.195 1.615 2.730 ;
        RECT  0.230 2.310 1.185 2.730 ;
        RECT  0.110 1.810 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.720 2.520 ;
        LAYER M1 ;
        RECT  6.330 1.000 6.390 1.260 ;
        RECT  6.210 1.000 6.330 1.900 ;
        RECT  5.700 1.780 6.210 1.900 ;
        RECT  5.580 0.395 5.700 1.900 ;
        RECT  5.495 0.395 5.580 0.565 ;
        RECT  4.945 1.780 5.580 1.900 ;
        RECT  5.320 1.260 5.440 1.520 ;
        RECT  4.460 1.260 5.320 1.380 ;
        RECT  4.940 1.550 4.945 1.900 ;
        RECT  4.825 1.500 4.940 1.900 ;
        RECT  4.680 1.500 4.825 1.620 ;
        RECT  4.310 2.020 4.570 2.190 ;
        RECT  4.420 0.640 4.515 0.760 ;
        RECT  4.450 1.260 4.460 1.805 ;
        RECT  4.420 1.260 4.450 1.900 ;
        RECT  4.300 0.640 4.420 1.900 ;
        RECT  3.780 2.020 4.310 2.140 ;
        RECT  4.255 0.640 4.300 0.760 ;
        RECT  4.190 1.780 4.300 1.900 ;
        RECT  4.020 0.650 4.055 1.460 ;
        RECT  3.935 0.650 4.020 1.870 ;
        RECT  3.900 1.340 3.935 1.870 ;
        RECT  3.090 1.340 3.900 1.460 ;
        RECT  3.660 1.590 3.780 2.140 ;
        RECT  2.940 1.590 3.660 1.710 ;
        RECT  3.130 1.865 3.250 2.190 ;
        RECT  2.380 1.865 3.130 1.985 ;
        RECT  2.975 0.620 3.095 1.220 ;
        RECT  2.275 0.620 2.975 0.740 ;
        RECT  2.940 1.100 2.975 1.220 ;
        RECT  2.820 1.100 2.940 1.710 ;
        RECT  2.485 0.860 2.855 0.980 ;
        RECT  2.380 0.860 2.485 1.565 ;
        RECT  2.365 0.860 2.380 2.010 ;
        RECT  2.260 1.445 2.365 2.010 ;
        RECT  2.140 0.620 2.275 0.780 ;
        RECT  0.470 1.890 2.260 2.010 ;
        RECT  2.135 0.980 2.195 1.240 ;
        RECT  2.135 0.660 2.140 0.780 ;
        RECT  2.015 0.660 2.135 1.760 ;
        RECT  0.710 1.640 2.015 1.760 ;
        RECT  1.775 0.660 1.895 1.520 ;
        RECT  1.240 0.660 1.775 0.780 ;
        RECT  1.000 1.400 1.775 1.520 ;
        RECT  0.880 1.000 1.000 1.520 ;
        RECT  0.710 1.000 0.880 1.120 ;
        RECT  0.590 0.760 0.710 1.120 ;
        RECT  0.590 1.240 0.710 1.760 ;
        RECT  0.430 0.760 0.590 0.880 ;
        RECT  0.350 1.000 0.470 2.010 ;
        RECT  0.310 0.620 0.430 0.880 ;
        RECT  0.190 1.000 0.350 1.120 ;
        RECT  0.190 0.380 0.330 0.500 ;
        RECT  0.070 0.380 0.190 1.120 ;
    END
END DFFRX1AD
MACRO DFFRX2AD
    CLASS CORE ;
    FOREIGN DFFRX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.085 0.920 5.255 1.095 ;
        RECT  4.805 0.920 5.085 1.040 ;
        RECT  4.685 0.400 4.805 1.040 ;
        RECT  3.890 0.400 4.685 0.520 ;
        RECT  3.770 0.400 3.890 0.700 ;
        RECT  3.600 0.580 3.770 0.700 ;
        RECT  3.410 0.580 3.600 1.130 ;
        RECT  3.340 0.380 3.410 1.130 ;
        RECT  3.290 0.380 3.340 0.700 ;
        RECT  2.170 0.380 3.290 0.500 ;
        RECT  2.050 0.380 2.170 0.540 ;
        RECT  1.050 0.420 2.050 0.540 ;
        RECT  0.875 0.420 1.050 0.880 ;
        END
        AntennaGateArea 0.112 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.025 0.390 6.195 1.660 ;
        RECT  5.950 0.860 6.025 1.355 ;
        END
        AntennaDiffArea 0.336 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.790 0.345 6.930 1.930 ;
        RECT  6.760 0.345 6.790 0.865 ;
        RECT  6.760 1.410 6.790 1.930 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 1.290 0.265 1.460 ;
        RECT  0.070 1.290 0.230 1.655 ;
        END
        AntennaGateArea 0.087 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.910 1.655 1.215 ;
        END
        AntennaGateArea 0.086 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.555 -0.210 7.000 0.210 ;
        RECT  6.385 -0.210 6.555 0.825 ;
        RECT  5.135 -0.210 6.385 0.210 ;
        RECT  4.965 -0.210 5.135 0.785 ;
        RECT  3.650 -0.210 4.965 0.210 ;
        RECT  3.530 -0.210 3.650 0.460 ;
        RECT  1.840 -0.210 3.530 0.210 ;
        RECT  1.580 -0.210 1.840 0.300 ;
        RECT  1.240 -0.210 1.580 0.210 ;
        RECT  0.980 -0.210 1.240 0.300 ;
        RECT  0.000 -0.210 0.980 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.555 2.310 7.000 2.730 ;
        RECT  6.385 2.055 6.555 2.730 ;
        RECT  5.875 2.310 6.385 2.730 ;
        RECT  5.705 2.020 5.875 2.730 ;
        RECT  5.205 2.310 5.705 2.730 ;
        RECT  4.945 2.210 5.205 2.730 ;
        RECT  3.590 2.310 4.945 2.730 ;
        RECT  3.420 1.830 3.590 2.730 ;
        RECT  3.010 2.310 3.420 2.730 ;
        RECT  2.750 2.130 3.010 2.730 ;
        RECT  1.805 2.310 2.750 2.730 ;
        RECT  1.635 2.165 1.805 2.730 ;
        RECT  1.245 2.310 1.635 2.730 ;
        RECT  1.075 2.145 1.245 2.730 ;
        RECT  0.230 2.310 1.075 2.730 ;
        RECT  0.110 1.810 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.570 1.000 6.670 1.260 ;
        RECT  6.450 1.000 6.570 1.900 ;
        RECT  5.830 1.780 6.450 1.900 ;
        RECT  5.710 0.585 5.830 1.900 ;
        RECT  5.575 0.585 5.710 0.755 ;
        RECT  5.060 1.780 5.710 1.900 ;
        RECT  5.470 1.010 5.590 1.530 ;
        RECT  4.420 1.260 5.470 1.380 ;
        RECT  4.940 1.500 5.060 1.900 ;
        RECT  4.800 1.500 4.940 1.620 ;
        RECT  4.620 2.060 4.690 2.180 ;
        RECT  4.430 2.020 4.620 2.180 ;
        RECT  4.420 1.780 4.570 1.900 ;
        RECT  4.420 0.640 4.565 0.760 ;
        RECT  3.830 2.020 4.430 2.140 ;
        RECT  4.300 0.640 4.420 1.900 ;
        RECT  4.010 0.660 4.130 1.870 ;
        RECT  3.950 1.340 4.010 1.870 ;
        RECT  3.090 1.340 3.950 1.460 ;
        RECT  3.710 1.590 3.830 2.140 ;
        RECT  2.940 1.590 3.710 1.710 ;
        RECT  3.130 1.830 3.250 2.190 ;
        RECT  2.700 1.830 3.130 1.950 ;
        RECT  2.975 0.620 3.095 1.220 ;
        RECT  2.460 0.620 2.975 0.740 ;
        RECT  2.940 1.100 2.975 1.220 ;
        RECT  2.820 1.100 2.940 1.710 ;
        RECT  2.700 0.860 2.840 0.980 ;
        RECT  2.580 0.860 2.700 1.950 ;
        RECT  2.430 1.830 2.580 1.950 ;
        RECT  2.340 0.620 2.460 1.520 ;
        RECT  2.380 1.675 2.430 1.950 ;
        RECT  2.260 1.675 2.380 2.010 ;
        RECT  2.015 0.665 2.340 0.835 ;
        RECT  1.865 1.400 2.340 1.520 ;
        RECT  0.505 1.890 2.260 2.010 ;
        RECT  1.895 0.990 2.200 1.250 ;
        RECT  1.775 0.660 1.895 1.250 ;
        RECT  1.745 1.400 1.865 1.760 ;
        RECT  1.290 0.660 1.775 0.780 ;
        RECT  0.745 1.640 1.745 1.760 ;
        RECT  1.290 1.400 1.470 1.520 ;
        RECT  1.170 0.660 1.290 1.520 ;
        RECT  0.745 1.000 1.170 1.120 ;
        RECT  0.625 0.790 0.745 1.120 ;
        RECT  0.625 1.250 0.745 1.760 ;
        RECT  0.430 0.790 0.625 0.910 ;
        RECT  0.385 1.030 0.505 2.010 ;
        RECT  0.310 0.650 0.430 0.910 ;
        RECT  0.190 1.030 0.385 1.150 ;
        RECT  0.190 0.380 0.350 0.500 ;
        RECT  0.070 0.380 0.190 1.150 ;
    END
END DFFRX2AD
MACRO DFFRX4AD
    CLASS CORE ;
    FOREIGN DFFRX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.290 0.920 5.460 1.140 ;
        RECT  5.010 0.920 5.290 1.040 ;
        RECT  4.890 0.380 5.010 1.040 ;
        RECT  4.060 0.380 4.890 0.500 ;
        RECT  3.940 0.380 4.060 0.940 ;
        RECT  3.850 0.820 3.940 0.940 ;
        RECT  3.580 0.820 3.850 1.130 ;
        RECT  3.460 0.380 3.580 1.130 ;
        RECT  2.275 0.380 3.460 0.500 ;
        RECT  2.155 0.380 2.275 0.635 ;
        RECT  1.050 0.515 2.155 0.635 ;
        RECT  0.910 0.515 1.050 0.865 ;
        RECT  0.875 0.695 0.910 0.865 ;
        END
        AntennaGateArea 0.157 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.505 0.390 6.675 1.660 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.380 0.985 7.490 1.515 ;
        RECT  7.240 0.345 7.380 1.930 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 1.290 0.265 1.460 ;
        RECT  0.070 1.290 0.230 1.655 ;
        END
        AntennaGateArea 0.104 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.865 1.890 1.215 ;
        RECT  1.575 1.000 1.750 1.215 ;
        END
        AntennaGateArea 0.127 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.730 -0.210 7.840 0.210 ;
        RECT  7.560 -0.210 7.730 0.865 ;
        RECT  7.035 -0.210 7.560 0.210 ;
        RECT  6.865 -0.210 7.035 0.825 ;
        RECT  6.315 -0.210 6.865 0.210 ;
        RECT  6.145 -0.210 6.315 0.820 ;
        RECT  5.340 -0.210 6.145 0.210 ;
        RECT  5.170 -0.210 5.340 0.705 ;
        RECT  3.820 -0.210 5.170 0.210 ;
        RECT  3.700 -0.210 3.820 0.700 ;
        RECT  1.990 -0.210 3.700 0.210 ;
        RECT  1.730 -0.210 1.990 0.395 ;
        RECT  1.210 -0.210 1.730 0.210 ;
        RECT  0.950 -0.210 1.210 0.390 ;
        RECT  0.000 -0.210 0.950 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.755 2.310 7.840 2.730 ;
        RECT  7.585 1.655 7.755 2.730 ;
        RECT  7.035 2.310 7.585 2.730 ;
        RECT  6.865 2.055 7.035 2.730 ;
        RECT  6.315 2.310 6.865 2.730 ;
        RECT  6.145 2.105 6.315 2.730 ;
        RECT  5.595 2.310 6.145 2.730 ;
        RECT  5.335 2.210 5.595 2.730 ;
        RECT  4.030 2.310 5.335 2.730 ;
        RECT  3.860 1.830 4.030 2.730 ;
        RECT  3.415 2.310 3.860 2.730 ;
        RECT  3.245 2.105 3.415 2.730 ;
        RECT  1.990 2.310 3.245 2.730 ;
        RECT  1.730 2.130 1.990 2.730 ;
        RECT  1.245 2.310 1.730 2.730 ;
        RECT  1.075 2.130 1.245 2.730 ;
        RECT  0.255 2.310 1.075 2.730 ;
        RECT  0.085 1.845 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.840 2.520 ;
        LAYER M1 ;
        RECT  7.050 1.000 7.100 1.260 ;
        RECT  6.930 1.000 7.050 1.900 ;
        RECT  6.345 1.780 6.930 1.900 ;
        RECT  6.225 0.940 6.345 1.900 ;
        RECT  5.950 0.940 6.225 1.060 ;
        RECT  5.500 1.780 6.225 1.900 ;
        RECT  5.885 1.185 6.055 1.615 ;
        RECT  5.830 0.535 5.950 1.060 ;
        RECT  4.895 1.260 5.885 1.380 ;
        RECT  5.780 0.535 5.830 0.705 ;
        RECT  5.380 1.500 5.500 1.900 ;
        RECT  5.240 1.500 5.380 1.620 ;
        RECT  5.060 2.060 5.130 2.180 ;
        RECT  4.870 2.020 5.060 2.180 ;
        RECT  4.750 1.260 4.895 1.870 ;
        RECT  4.270 2.020 4.870 2.140 ;
        RECT  4.745 0.640 4.750 1.870 ;
        RECT  4.630 0.640 4.745 1.380 ;
        RECT  4.490 0.640 4.630 0.760 ;
        RECT  4.390 1.340 4.510 1.870 ;
        RECT  4.300 1.340 4.390 1.460 ;
        RECT  4.180 0.660 4.300 1.460 ;
        RECT  4.150 1.590 4.270 2.140 ;
        RECT  3.350 1.340 4.180 1.460 ;
        RECT  3.230 1.590 4.150 1.710 ;
        RECT  3.615 1.830 3.735 2.190 ;
        RECT  2.835 1.830 3.615 1.950 ;
        RECT  3.230 0.620 3.335 1.220 ;
        RECT  3.215 0.620 3.230 1.710 ;
        RECT  2.580 0.620 3.215 0.740 ;
        RECT  3.110 1.100 3.215 1.710 ;
        RECT  2.820 0.860 3.080 0.980 ;
        RECT  2.820 1.675 2.835 1.950 ;
        RECT  2.735 0.860 2.820 1.950 ;
        RECT  2.700 0.860 2.735 2.010 ;
        RECT  2.615 1.675 2.700 2.010 ;
        RECT  0.505 1.890 2.615 2.010 ;
        RECT  2.470 0.620 2.580 1.520 ;
        RECT  2.460 0.620 2.470 1.760 ;
        RECT  2.090 0.755 2.460 0.875 ;
        RECT  2.350 1.400 2.460 1.760 ;
        RECT  0.745 1.640 2.350 1.760 ;
        RECT  2.060 1.045 2.230 1.520 ;
        RECT  1.440 1.400 2.060 1.520 ;
        RECT  1.440 0.755 1.580 0.875 ;
        RECT  1.320 0.755 1.440 1.520 ;
        RECT  0.745 1.000 1.320 1.120 ;
        RECT  0.625 0.790 0.745 1.120 ;
        RECT  0.625 1.250 0.745 1.760 ;
        RECT  0.430 0.790 0.625 0.910 ;
        RECT  0.385 1.030 0.505 2.010 ;
        RECT  0.310 0.650 0.430 0.910 ;
        RECT  0.190 1.030 0.385 1.150 ;
        RECT  0.190 0.380 0.350 0.500 ;
        RECT  0.070 0.380 0.190 1.150 ;
    END
END DFFRX4AD
MACRO DFFRXLAD
    CLASS CORE ;
    FOREIGN DFFRXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 0.400 5.160 1.140 ;
        RECT  3.815 0.400 5.040 0.520 ;
        RECT  3.695 0.400 3.815 0.760 ;
        RECT  3.590 0.640 3.695 0.760 ;
        RECT  3.470 0.640 3.590 1.220 ;
        RECT  3.335 0.640 3.470 0.760 ;
        RECT  3.215 0.380 3.335 0.760 ;
        RECT  2.020 0.380 3.215 0.500 ;
        RECT  1.900 0.380 2.020 0.540 ;
        RECT  1.050 0.420 1.900 0.540 ;
        RECT  0.870 0.420 1.050 0.880 ;
        END
        AntennaGateArea 0.102 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.940 0.585 6.090 0.865 ;
        RECT  5.820 0.585 5.940 1.590 ;
        END
        AntennaDiffArea 0.132 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.510 0.735 6.650 1.690 ;
        RECT  6.465 0.735 6.510 0.905 ;
        RECT  6.485 1.410 6.510 1.690 ;
        END
        AntennaDiffArea 0.143 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.240 0.230 1.655 ;
        END
        AntennaGateArea 0.067 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.910 1.655 1.060 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.290 -0.210 6.720 0.210 ;
        RECT  6.030 -0.210 6.290 0.430 ;
        RECT  5.060 -0.210 6.030 0.210 ;
        RECT  4.800 -0.210 5.060 0.280 ;
        RECT  3.575 -0.210 4.800 0.210 ;
        RECT  3.455 -0.210 3.575 0.475 ;
        RECT  1.780 -0.210 3.455 0.210 ;
        RECT  1.520 -0.210 1.780 0.300 ;
        RECT  1.240 -0.210 1.520 0.210 ;
        RECT  0.980 -0.210 1.240 0.300 ;
        RECT  0.000 -0.210 0.980 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.255 2.310 6.720 2.730 ;
        RECT  6.085 2.020 6.255 2.730 ;
        RECT  5.755 2.310 6.085 2.730 ;
        RECT  5.585 2.020 5.755 2.730 ;
        RECT  5.035 2.310 5.585 2.730 ;
        RECT  4.775 2.210 5.035 2.730 ;
        RECT  3.540 2.310 4.775 2.730 ;
        RECT  3.370 1.830 3.540 2.730 ;
        RECT  3.010 2.310 3.370 2.730 ;
        RECT  2.750 2.105 3.010 2.730 ;
        RECT  1.715 2.310 2.750 2.730 ;
        RECT  1.545 2.165 1.715 2.730 ;
        RECT  1.245 2.310 1.545 2.730 ;
        RECT  1.075 2.130 1.245 2.730 ;
        RECT  0.230 2.310 1.075 2.730 ;
        RECT  0.110 1.810 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.720 2.520 ;
        LAYER M1 ;
        RECT  6.330 1.000 6.390 1.260 ;
        RECT  6.210 1.000 6.330 1.900 ;
        RECT  5.700 1.780 6.210 1.900 ;
        RECT  5.580 0.395 5.700 1.900 ;
        RECT  5.495 0.395 5.580 0.565 ;
        RECT  4.945 1.780 5.580 1.900 ;
        RECT  5.320 1.260 5.440 1.520 ;
        RECT  4.460 1.260 5.320 1.380 ;
        RECT  4.940 1.550 4.945 1.900 ;
        RECT  4.825 1.500 4.940 1.900 ;
        RECT  4.680 1.500 4.825 1.620 ;
        RECT  4.310 2.020 4.570 2.190 ;
        RECT  4.420 0.640 4.515 0.760 ;
        RECT  4.450 1.260 4.460 1.805 ;
        RECT  4.420 1.260 4.450 1.900 ;
        RECT  4.300 0.640 4.420 1.900 ;
        RECT  3.780 2.020 4.310 2.140 ;
        RECT  4.255 0.640 4.300 0.760 ;
        RECT  4.190 1.780 4.300 1.900 ;
        RECT  4.020 0.650 4.055 1.460 ;
        RECT  3.935 0.650 4.020 1.870 ;
        RECT  3.900 1.340 3.935 1.870 ;
        RECT  3.090 1.340 3.900 1.460 ;
        RECT  3.660 1.590 3.780 2.140 ;
        RECT  2.940 1.590 3.660 1.710 ;
        RECT  3.130 1.865 3.250 2.190 ;
        RECT  2.380 1.865 3.130 1.985 ;
        RECT  2.975 0.620 3.095 1.220 ;
        RECT  2.275 0.620 2.975 0.740 ;
        RECT  2.940 1.100 2.975 1.220 ;
        RECT  2.820 1.100 2.940 1.710 ;
        RECT  2.485 0.860 2.855 0.980 ;
        RECT  2.380 0.860 2.485 1.565 ;
        RECT  2.365 0.860 2.380 2.010 ;
        RECT  2.260 1.445 2.365 2.010 ;
        RECT  2.140 0.620 2.275 0.780 ;
        RECT  0.470 1.890 2.260 2.010 ;
        RECT  2.135 0.980 2.195 1.240 ;
        RECT  2.135 0.660 2.140 0.780 ;
        RECT  2.015 0.660 2.135 1.760 ;
        RECT  0.710 1.640 2.015 1.760 ;
        RECT  1.775 0.660 1.895 1.520 ;
        RECT  1.240 0.660 1.775 0.780 ;
        RECT  0.950 1.400 1.775 1.520 ;
        RECT  0.830 1.000 0.950 1.520 ;
        RECT  0.710 1.000 0.830 1.120 ;
        RECT  0.590 0.760 0.710 1.120 ;
        RECT  0.590 1.240 0.710 1.760 ;
        RECT  0.430 0.760 0.590 0.880 ;
        RECT  0.350 1.000 0.470 2.010 ;
        RECT  0.310 0.620 0.430 0.880 ;
        RECT  0.190 1.000 0.350 1.120 ;
        RECT  0.190 0.380 0.330 0.500 ;
        RECT  0.070 0.380 0.190 1.120 ;
    END
END DFFRXLAD
MACRO DFFSHQX1AD
    CLASS CORE ;
    FOREIGN DFFSHQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 0.870 3.040 1.375 ;
        RECT  2.660 0.960 2.870 1.220 ;
        END
        AntennaGateArea 0.109 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.610 0.600 7.770 1.930 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 0.865 1.990 1.185 ;
        RECT  1.750 0.865 1.890 1.370 ;
        END
        AntennaGateArea 0.048 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.000 0.530 1.375 ;
        END
        AntennaGateArea 0.118 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.375 -0.210 7.840 0.210 ;
        RECT  7.205 -0.210 7.375 0.335 ;
        RECT  6.545 -0.210 7.205 0.210 ;
        RECT  6.285 -0.210 6.545 0.330 ;
        RECT  4.700 -0.210 6.285 0.210 ;
        RECT  4.530 -0.210 4.700 0.260 ;
        RECT  2.935 -0.210 4.530 0.210 ;
        RECT  2.675 -0.210 2.935 0.260 ;
        RECT  1.915 -0.210 2.675 0.210 ;
        RECT  1.745 -0.210 1.915 0.260 ;
        RECT  1.165 -0.210 1.745 0.210 ;
        RECT  0.995 -0.210 1.165 0.375 ;
        RECT  0.635 -0.210 0.995 0.210 ;
        RECT  0.465 -0.210 0.635 0.375 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.330 2.310 7.840 2.730 ;
        RECT  6.890 1.965 7.330 2.730 ;
        RECT  5.170 2.310 6.890 2.730 ;
        RECT  5.000 1.925 5.170 2.730 ;
        RECT  4.035 2.310 5.000 2.730 ;
        RECT  3.915 2.145 4.035 2.730 ;
        RECT  2.840 2.310 3.915 2.730 ;
        RECT  2.670 2.145 2.840 2.730 ;
        RECT  1.870 2.310 2.670 2.730 ;
        RECT  1.700 2.145 1.870 2.730 ;
        RECT  0.530 2.310 1.700 2.730 ;
        RECT  0.410 1.780 0.530 2.730 ;
        RECT  0.000 2.310 0.410 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.840 2.520 ;
        LAYER M1 ;
        RECT  7.245 0.455 7.365 1.840 ;
        RECT  6.880 0.455 7.245 0.575 ;
        RECT  6.715 1.720 7.245 1.840 ;
        RECT  6.855 0.695 7.025 1.545 ;
        RECT  6.710 0.355 6.880 0.575 ;
        RECT  6.595 1.070 6.855 1.240 ;
        RECT  6.595 1.720 6.715 2.045 ;
        RECT  5.725 0.455 6.710 0.575 ;
        RECT  6.475 0.755 6.685 0.875 ;
        RECT  5.765 1.925 6.595 2.045 ;
        RECT  6.355 0.755 6.475 1.805 ;
        RECT  4.755 1.685 6.355 1.805 ;
        RECT  6.055 0.925 6.175 1.565 ;
        RECT  5.485 0.925 6.055 1.045 ;
        RECT  5.605 0.455 5.725 0.720 ;
        RECT  5.205 1.405 5.645 1.565 ;
        RECT  5.365 0.380 5.485 1.045 ;
        RECT  4.115 0.380 5.365 0.500 ;
        RECT  5.085 0.670 5.205 1.565 ;
        RECT  4.875 1.375 5.085 1.565 ;
        RECT  4.845 0.620 4.965 1.255 ;
        RECT  2.490 0.620 4.845 0.740 ;
        RECT  4.755 1.135 4.845 1.255 ;
        RECT  4.635 1.135 4.755 1.805 ;
        RECT  3.965 0.895 4.725 1.015 ;
        RECT  4.445 2.020 4.705 2.190 ;
        RECT  4.395 1.490 4.515 1.900 ;
        RECT  4.275 2.020 4.445 2.140 ;
        RECT  3.825 1.490 4.395 1.610 ;
        RECT  4.155 1.905 4.275 2.140 ;
        RECT  3.375 1.905 4.155 2.025 ;
        RECT  3.855 0.335 4.115 0.500 ;
        RECT  3.825 0.860 3.965 1.015 ;
        RECT  1.550 0.380 3.855 0.500 ;
        RECT  3.705 0.860 3.825 1.610 ;
        RECT  3.625 1.490 3.705 1.610 ;
        RECT  3.505 1.490 3.625 1.750 ;
        RECT  3.375 0.935 3.420 1.055 ;
        RECT  3.255 0.935 3.375 2.025 ;
        RECT  3.160 0.935 3.255 1.055 ;
        RECT  1.160 1.905 3.255 2.025 ;
        RECT  2.930 1.615 3.100 1.785 ;
        RECT  2.250 1.665 2.930 1.785 ;
        RECT  2.490 1.375 2.545 1.545 ;
        RECT  2.370 0.620 2.490 1.545 ;
        RECT  2.130 0.625 2.250 1.785 ;
        RECT  1.990 0.625 2.130 0.745 ;
        RECT  2.035 1.415 2.130 1.585 ;
        RECT  1.430 0.335 1.550 1.520 ;
        RECT  1.010 1.400 1.430 1.520 ;
        RECT  1.190 0.495 1.310 1.195 ;
        RECT  0.230 0.495 1.190 0.615 ;
        RECT  1.040 1.670 1.160 2.025 ;
        RECT  0.770 1.670 1.040 1.790 ;
        RECT  0.890 1.020 1.010 1.520 ;
        RECT  0.770 0.760 0.980 0.880 ;
        RECT  0.650 0.760 0.770 1.790 ;
        RECT  0.110 0.495 0.230 1.600 ;
    END
END DFFSHQX1AD
MACRO DFFSHQX2AD
    CLASS CORE ;
    FOREIGN DFFSHQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 0.870 3.040 1.375 ;
        RECT  2.660 0.980 2.870 1.240 ;
        END
        AntennaGateArea 0.137 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.610 0.600 7.770 2.190 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 0.865 1.990 1.185 ;
        RECT  1.750 0.865 1.890 1.370 ;
        END
        AntennaGateArea 0.048 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.000 0.530 1.375 ;
        END
        AntennaGateArea 0.121 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.325 -0.210 7.840 0.210 ;
        RECT  7.155 -0.210 7.325 0.335 ;
        RECT  6.545 -0.210 7.155 0.210 ;
        RECT  6.285 -0.210 6.545 0.330 ;
        RECT  4.700 -0.210 6.285 0.210 ;
        RECT  4.530 -0.210 4.700 0.260 ;
        RECT  2.935 -0.210 4.530 0.210 ;
        RECT  2.675 -0.210 2.935 0.260 ;
        RECT  1.915 -0.210 2.675 0.210 ;
        RECT  1.745 -0.210 1.915 0.260 ;
        RECT  1.165 -0.210 1.745 0.210 ;
        RECT  0.995 -0.210 1.165 0.375 ;
        RECT  0.635 -0.210 0.995 0.210 ;
        RECT  0.465 -0.210 0.635 0.375 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.325 2.310 7.840 2.730 ;
        RECT  6.895 1.960 7.325 2.730 ;
        RECT  5.170 2.310 6.895 2.730 ;
        RECT  5.000 1.925 5.170 2.730 ;
        RECT  4.280 2.310 5.000 2.730 ;
        RECT  4.110 2.265 4.280 2.730 ;
        RECT  2.840 2.310 4.110 2.730 ;
        RECT  2.670 2.260 2.840 2.730 ;
        RECT  1.870 2.310 2.670 2.730 ;
        RECT  1.700 2.260 1.870 2.730 ;
        RECT  0.530 2.310 1.700 2.730 ;
        RECT  0.410 1.780 0.530 2.730 ;
        RECT  0.000 2.310 0.410 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.840 2.520 ;
        LAYER M1 ;
        RECT  7.245 0.455 7.365 1.840 ;
        RECT  6.880 0.455 7.245 0.575 ;
        RECT  6.715 1.720 7.245 1.840 ;
        RECT  6.855 0.735 7.025 1.545 ;
        RECT  6.710 0.355 6.880 0.575 ;
        RECT  6.595 1.070 6.855 1.240 ;
        RECT  6.595 1.720 6.715 2.045 ;
        RECT  5.725 0.455 6.710 0.575 ;
        RECT  6.475 0.755 6.685 0.875 ;
        RECT  5.765 1.925 6.595 2.045 ;
        RECT  6.355 0.755 6.475 1.805 ;
        RECT  4.755 1.685 6.355 1.805 ;
        RECT  6.055 0.925 6.175 1.565 ;
        RECT  5.485 0.925 6.055 1.045 ;
        RECT  5.605 0.455 5.725 0.720 ;
        RECT  5.205 1.405 5.645 1.545 ;
        RECT  5.365 0.380 5.485 1.045 ;
        RECT  4.115 0.380 5.365 0.500 ;
        RECT  5.085 0.620 5.205 1.545 ;
        RECT  4.875 1.375 5.085 1.545 ;
        RECT  4.845 0.620 4.965 1.255 ;
        RECT  2.490 0.620 4.845 0.740 ;
        RECT  4.755 1.135 4.845 1.255 ;
        RECT  4.635 1.135 4.755 1.805 ;
        RECT  3.965 0.895 4.725 1.015 ;
        RECT  4.445 2.020 4.705 2.190 ;
        RECT  4.395 1.490 4.515 1.900 ;
        RECT  3.385 2.020 4.445 2.140 ;
        RECT  3.825 1.490 4.395 1.610 ;
        RECT  3.855 0.335 4.115 0.500 ;
        RECT  3.825 0.860 3.965 1.015 ;
        RECT  1.550 0.380 3.855 0.500 ;
        RECT  3.705 0.860 3.825 1.610 ;
        RECT  3.625 1.490 3.705 1.610 ;
        RECT  3.505 1.490 3.625 1.785 ;
        RECT  3.385 1.045 3.420 1.165 ;
        RECT  3.265 1.045 3.385 2.140 ;
        RECT  3.160 1.045 3.265 1.165 ;
        RECT  1.160 2.020 3.265 2.140 ;
        RECT  2.250 1.780 3.145 1.900 ;
        RECT  2.490 1.375 2.545 1.545 ;
        RECT  2.370 0.620 2.490 1.545 ;
        RECT  2.130 0.625 2.250 1.900 ;
        RECT  1.990 0.625 2.130 0.745 ;
        RECT  2.035 1.415 2.130 1.585 ;
        RECT  1.430 0.330 1.550 1.520 ;
        RECT  1.010 1.400 1.430 1.520 ;
        RECT  1.190 0.495 1.310 1.195 ;
        RECT  0.230 0.495 1.190 0.615 ;
        RECT  1.040 1.670 1.160 2.140 ;
        RECT  0.770 1.670 1.040 1.790 ;
        RECT  0.890 1.020 1.010 1.520 ;
        RECT  0.770 0.760 0.980 0.880 ;
        RECT  0.650 0.760 0.770 1.790 ;
        RECT  0.110 0.495 0.230 1.600 ;
    END
END DFFSHQX2AD
MACRO DFFSHQX4AD
    CLASS CORE ;
    FOREIGN DFFSHQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 0.960 3.010 1.375 ;
        END
        AntennaGateArea 0.156 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.795 1.005 8.890 1.515 ;
        RECT  8.625 0.415 8.795 2.170 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 0.865 1.950 1.060 ;
        RECT  1.470 0.865 1.890 1.095 ;
        END
        AntennaGateArea 0.079 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.325 0.870 0.490 1.445 ;
        END
        AntennaGateArea 0.192 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.155 -0.210 9.240 0.210 ;
        RECT  8.985 -0.210 9.155 0.845 ;
        RECT  8.365 -0.210 8.985 0.210 ;
        RECT  8.195 -0.210 8.365 0.270 ;
        RECT  7.455 -0.210 8.195 0.210 ;
        RECT  7.285 -0.210 7.455 0.325 ;
        RECT  5.780 -0.210 7.285 0.210 ;
        RECT  5.520 -0.210 5.780 0.630 ;
        RECT  4.880 -0.210 5.520 0.210 ;
        RECT  4.620 -0.210 4.880 0.500 ;
        RECT  2.930 -0.210 4.620 0.210 ;
        RECT  2.760 -0.210 2.930 0.260 ;
        RECT  1.815 -0.210 2.760 0.210 ;
        RECT  1.555 -0.210 1.815 0.230 ;
        RECT  0.635 -0.210 1.555 0.210 ;
        RECT  0.465 -0.210 0.635 0.255 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.155 2.310 9.240 2.730 ;
        RECT  8.985 1.635 9.155 2.730 ;
        RECT  8.435 2.310 8.985 2.730 ;
        RECT  8.005 1.960 8.435 2.730 ;
        RECT  6.105 2.310 8.005 2.730 ;
        RECT  5.935 1.910 6.105 2.730 ;
        RECT  5.295 2.310 5.935 2.730 ;
        RECT  5.125 1.910 5.295 2.730 ;
        RECT  4.355 2.310 5.125 2.730 ;
        RECT  4.095 2.260 4.355 2.730 ;
        RECT  2.825 2.310 4.095 2.730 ;
        RECT  2.655 2.260 2.825 2.730 ;
        RECT  1.880 2.310 2.655 2.730 ;
        RECT  1.620 2.260 1.880 2.730 ;
        RECT  0.575 2.310 1.620 2.730 ;
        RECT  0.405 2.075 0.575 2.730 ;
        RECT  0.000 2.310 0.405 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.240 2.520 ;
        LAYER M1 ;
        RECT  8.345 0.445 8.465 1.840 ;
        RECT  6.825 0.445 8.345 0.565 ;
        RECT  7.885 1.720 8.345 1.840 ;
        RECT  7.980 0.690 8.100 1.590 ;
        RECT  7.890 1.025 7.980 1.285 ;
        RECT  7.765 1.720 7.885 2.055 ;
        RECT  7.630 0.755 7.770 0.875 ;
        RECT  6.230 1.935 7.765 2.055 ;
        RECT  7.510 0.755 7.630 1.790 ;
        RECT  4.840 1.670 7.510 1.790 ;
        RECT  7.210 1.040 7.330 1.525 ;
        RECT  6.360 1.040 7.210 1.160 ;
        RECT  5.350 1.430 6.850 1.550 ;
        RECT  6.655 0.380 6.825 0.565 ;
        RECT  6.105 0.380 6.655 0.500 ;
        RECT  6.250 0.620 6.510 0.870 ;
        RECT  6.100 0.990 6.360 1.160 ;
        RECT  5.350 0.750 6.250 0.870 ;
        RECT  5.935 0.380 6.105 0.630 ;
        RECT  5.230 0.540 5.350 1.550 ;
        RECT  4.960 1.390 5.230 1.550 ;
        RECT  4.990 0.620 5.110 1.270 ;
        RECT  2.440 0.620 4.990 0.740 ;
        RECT  4.840 1.150 4.990 1.270 ;
        RECT  4.600 0.860 4.860 1.030 ;
        RECT  4.720 1.150 4.840 1.790 ;
        RECT  4.565 2.020 4.825 2.190 ;
        RECT  3.920 0.860 4.600 0.980 ;
        RECT  4.430 1.575 4.600 1.855 ;
        RECT  3.415 2.020 4.565 2.140 ;
        RECT  3.920 1.575 4.430 1.695 ;
        RECT  3.960 0.330 4.220 0.500 ;
        RECT  1.800 0.380 3.960 0.500 ;
        RECT  3.800 0.860 3.920 1.695 ;
        RECT  3.655 1.510 3.800 1.695 ;
        RECT  3.535 1.510 3.655 1.770 ;
        RECT  3.415 1.030 3.580 1.150 ;
        RECT  3.295 1.030 3.415 2.140 ;
        RECT  1.160 2.020 3.295 2.140 ;
        RECT  2.195 1.780 3.130 1.900 ;
        RECT  2.320 0.620 2.440 1.590 ;
        RECT  2.075 0.620 2.195 1.900 ;
        RECT  1.935 0.620 2.075 0.740 ;
        RECT  1.980 1.200 2.075 1.720 ;
        RECT  1.680 0.380 1.800 0.740 ;
        RECT  1.150 0.620 1.680 0.740 ;
        RECT  1.210 0.330 1.470 0.500 ;
        RECT  1.285 1.220 1.455 1.545 ;
        RECT  1.150 1.220 1.285 1.340 ;
        RECT  0.670 0.380 1.210 0.500 ;
        RECT  1.040 1.670 1.160 2.190 ;
        RECT  1.030 0.620 1.150 1.340 ;
        RECT  0.730 1.670 1.040 1.790 ;
        RECT  0.850 1.220 1.030 1.340 ;
        RECT  0.790 0.620 0.910 1.000 ;
        RECT  0.730 0.875 0.790 1.000 ;
        RECT  0.610 0.875 0.730 1.790 ;
        RECT  0.550 0.380 0.670 0.750 ;
        RECT  0.255 0.630 0.550 0.750 ;
        RECT  0.205 0.580 0.255 0.750 ;
        RECT  0.205 1.560 0.255 1.730 ;
        RECT  0.085 0.580 0.205 1.730 ;
    END
END DFFSHQX4AD
MACRO DFFSHQX8AD
    CLASS CORE ;
    FOREIGN DFFSHQX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.065 0.960 3.455 1.375 ;
        END
        AntennaGateArea 0.166 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.905 0.370 10.075 2.170 ;
        RECT  9.355 1.005 9.905 1.515 ;
        RECT  9.170 0.370 9.355 2.170 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 0.865 2.235 1.250 ;
        END
        AntennaGateArea 0.143 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.025 0.790 1.375 ;
        END
        AntennaGateArea 0.29 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.435 -0.210 10.640 0.210 ;
        RECT  10.265 -0.210 10.435 0.800 ;
        RECT  9.715 -0.210 10.265 0.210 ;
        RECT  9.545 -0.210 9.715 0.800 ;
        RECT  8.995 -0.210 9.545 0.210 ;
        RECT  8.825 -0.210 8.995 0.800 ;
        RECT  7.765 -0.210 8.825 0.210 ;
        RECT  7.595 -0.210 7.765 0.325 ;
        RECT  6.060 -0.210 7.595 0.210 ;
        RECT  5.800 -0.210 6.060 0.630 ;
        RECT  5.160 -0.210 5.800 0.210 ;
        RECT  4.900 -0.210 5.160 0.500 ;
        RECT  3.295 -0.210 4.900 0.210 ;
        RECT  3.035 -0.210 3.295 0.260 ;
        RECT  1.855 -0.210 3.035 0.210 ;
        RECT  1.735 -0.210 1.855 0.500 ;
        RECT  0.790 -0.210 1.735 0.210 ;
        RECT  0.530 -0.210 0.790 0.260 ;
        RECT  0.000 -0.210 0.530 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.435 2.310 10.640 2.730 ;
        RECT  10.265 1.480 10.435 2.730 ;
        RECT  9.715 2.310 10.265 2.730 ;
        RECT  9.545 1.740 9.715 2.730 ;
        RECT  8.890 2.310 9.545 2.730 ;
        RECT  8.460 1.960 8.890 2.730 ;
        RECT  6.410 2.310 8.460 2.730 ;
        RECT  6.240 1.910 6.410 2.730 ;
        RECT  5.600 2.310 6.240 2.730 ;
        RECT  5.430 1.910 5.600 2.730 ;
        RECT  4.635 2.310 5.430 2.730 ;
        RECT  4.375 2.190 4.635 2.730 ;
        RECT  3.105 2.310 4.375 2.730 ;
        RECT  2.935 2.260 3.105 2.730 ;
        RECT  2.095 2.310 2.935 2.730 ;
        RECT  1.835 2.260 2.095 2.730 ;
        RECT  0.720 2.310 1.835 2.730 ;
        RECT  0.550 1.495 0.720 2.730 ;
        RECT  0.000 2.310 0.550 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.640 2.520 ;
        LAYER M1 ;
        RECT  8.760 0.990 9.020 1.250 ;
        RECT  8.705 0.990 8.760 1.840 ;
        RECT  8.640 0.445 8.705 1.840 ;
        RECT  8.585 0.445 8.640 1.250 ;
        RECT  8.230 1.720 8.640 1.840 ;
        RECT  7.105 0.445 8.585 0.565 ;
        RECT  8.465 1.375 8.520 1.545 ;
        RECT  8.345 0.690 8.465 1.545 ;
        RECT  8.305 1.070 8.345 1.545 ;
        RECT  8.130 1.070 8.305 1.235 ;
        RECT  8.110 1.720 8.230 2.055 ;
        RECT  7.990 0.790 8.130 0.910 ;
        RECT  6.535 1.935 8.110 2.055 ;
        RECT  7.870 0.790 7.990 1.790 ;
        RECT  5.145 1.670 7.870 1.790 ;
        RECT  7.560 1.040 7.680 1.550 ;
        RECT  6.670 1.040 7.560 1.160 ;
        RECT  5.630 1.430 7.160 1.550 ;
        RECT  6.935 0.380 7.105 0.565 ;
        RECT  6.385 0.380 6.935 0.500 ;
        RECT  6.530 0.620 6.790 0.870 ;
        RECT  6.410 0.990 6.670 1.160 ;
        RECT  5.630 0.750 6.530 0.870 ;
        RECT  6.215 0.380 6.385 0.630 ;
        RECT  5.510 0.540 5.630 1.550 ;
        RECT  5.265 1.430 5.510 1.550 ;
        RECT  5.270 0.620 5.390 1.310 ;
        RECT  2.745 0.620 5.270 0.740 ;
        RECT  5.145 1.190 5.270 1.310 ;
        RECT  5.025 1.190 5.145 1.790 ;
        RECT  4.880 0.860 5.140 1.070 ;
        RECT  4.845 1.950 5.105 2.190 ;
        RECT  4.645 1.575 4.905 1.830 ;
        RECT  4.200 0.860 4.880 0.980 ;
        RECT  3.695 1.950 4.845 2.070 ;
        RECT  4.200 1.575 4.645 1.695 ;
        RECT  4.240 0.330 4.500 0.500 ;
        RECT  2.095 0.380 4.240 0.500 ;
        RECT  4.080 0.860 4.200 1.695 ;
        RECT  3.935 1.510 4.080 1.695 ;
        RECT  3.815 1.510 3.935 1.770 ;
        RECT  3.695 1.030 3.860 1.150 ;
        RECT  3.575 1.030 3.695 2.140 ;
        RECT  1.305 2.020 3.575 2.140 ;
        RECT  2.475 1.780 3.410 1.900 ;
        RECT  2.625 0.620 2.745 1.585 ;
        RECT  2.355 0.625 2.475 1.900 ;
        RECT  2.215 0.625 2.355 0.745 ;
        RECT  2.260 1.470 2.355 1.900 ;
        RECT  1.975 0.380 2.095 0.740 ;
        RECT  1.670 0.620 1.975 0.740 ;
        RECT  1.500 0.620 1.670 1.900 ;
        RECT  1.305 0.620 1.500 0.740 ;
        RECT  1.265 1.055 1.500 1.315 ;
        RECT  1.100 0.330 1.360 0.500 ;
        RECT  1.185 1.485 1.305 2.140 ;
        RECT  1.100 1.485 1.185 1.605 ;
        RECT  0.360 0.380 1.100 0.500 ;
        RECT  0.980 0.620 1.100 1.605 ;
        RECT  0.190 0.380 0.360 0.810 ;
        RECT  0.190 1.495 0.360 1.925 ;
        RECT  0.070 0.595 0.190 1.710 ;
    END
END DFFSHQX8AD
MACRO DFFSQX1AD
    CLASS CORE ;
    FOREIGN DFFSQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.495 1.275 4.755 1.655 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.495 5.810 2.070 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 1.020 0.490 1.395 ;
        END
        AntennaGateArea 0.048 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.470 0.865 2.730 1.095 ;
        RECT  2.350 0.865 2.470 1.270 ;
        END
        AntennaGateArea 0.089 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.435 -0.210 5.880 0.210 ;
        RECT  5.265 -0.210 5.435 0.670 ;
        RECT  4.685 -0.210 5.265 0.210 ;
        RECT  4.515 -0.210 4.685 0.715 ;
        RECT  2.270 -0.210 4.515 0.210 ;
        RECT  2.010 -0.210 2.270 0.300 ;
        RECT  1.430 -0.210 2.010 0.210 ;
        RECT  1.170 -0.210 1.430 0.415 ;
        RECT  0.265 -0.210 1.170 0.210 ;
        RECT  0.095 -0.210 0.265 0.440 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.425 2.310 5.880 2.730 ;
        RECT  5.165 2.015 5.425 2.730 ;
        RECT  4.440 2.310 5.165 2.730 ;
        RECT  4.270 2.055 4.440 2.730 ;
        RECT  3.400 2.310 4.270 2.730 ;
        RECT  3.140 2.020 3.400 2.730 ;
        RECT  2.610 2.310 3.140 2.730 ;
        RECT  2.350 1.965 2.610 2.730 ;
        RECT  1.285 2.310 2.350 2.730 ;
        RECT  1.165 1.995 1.285 2.730 ;
        RECT  0.265 2.310 1.165 2.730 ;
        RECT  0.095 1.650 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.880 2.520 ;
        LAYER M1 ;
        RECT  5.410 0.790 5.530 1.895 ;
        RECT  5.085 0.790 5.410 0.910 ;
        RECT  4.900 1.775 5.410 1.895 ;
        RECT  4.915 0.665 5.085 0.910 ;
        RECT  4.905 1.030 5.065 1.595 ;
        RECT  3.825 1.030 4.905 1.150 ;
        RECT  4.730 1.775 4.900 2.105 ;
        RECT  4.355 1.775 4.730 1.895 ;
        RECT  4.230 1.315 4.355 1.895 ;
        RECT  4.155 0.380 4.325 0.725 ;
        RECT  4.095 1.315 4.230 1.435 ;
        RECT  2.590 0.380 4.155 0.500 ;
        RECT  3.925 1.780 4.045 2.140 ;
        RECT  3.525 1.780 3.925 1.900 ;
        RECT  3.705 0.620 3.825 1.660 ;
        RECT  3.435 0.620 3.705 0.740 ;
        RECT  3.645 1.390 3.705 1.660 ;
        RECT  3.525 0.860 3.550 1.120 ;
        RECT  3.405 0.860 3.525 1.900 ;
        RECT  1.770 1.725 3.405 1.845 ;
        RECT  3.165 0.620 3.285 1.575 ;
        RECT  2.470 0.620 3.165 0.740 ;
        RECT  2.830 1.455 3.165 1.575 ;
        RECT  2.900 1.070 3.020 1.335 ;
        RECT  2.710 1.215 2.900 1.335 ;
        RECT  2.590 1.215 2.710 1.605 ;
        RECT  2.230 1.485 2.590 1.605 ;
        RECT  2.350 0.420 2.470 0.740 ;
        RECT  1.990 0.420 2.350 0.540 ;
        RECT  2.110 0.660 2.230 1.605 ;
        RECT  2.005 1.145 2.110 1.605 ;
        RECT  1.525 2.020 2.030 2.140 ;
        RECT  1.440 1.145 2.005 1.265 ;
        RECT  1.870 0.420 1.990 1.025 ;
        RECT  1.295 0.905 1.870 1.025 ;
        RECT  1.650 1.385 1.770 1.845 ;
        RECT  1.630 0.525 1.750 0.785 ;
        RECT  1.055 1.385 1.650 1.505 ;
        RECT  1.055 0.665 1.630 0.785 ;
        RECT  1.405 1.625 1.525 2.140 ;
        RECT  0.740 1.625 1.405 1.745 ;
        RECT  1.175 0.905 1.295 1.225 ;
        RECT  0.935 0.665 1.055 1.505 ;
        RECT  0.860 1.045 0.935 1.505 ;
        RECT  0.740 0.655 0.815 0.915 ;
        RECT  0.620 0.655 0.740 1.745 ;
    END
END DFFSQX1AD
MACRO DFFSQX2AD
    CLASS CORE ;
    FOREIGN DFFSQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.495 1.275 4.755 1.655 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.650 0.380 5.810 1.985 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 1.020 0.490 1.395 ;
        END
        AntennaGateArea 0.048 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.470 0.865 2.730 1.095 ;
        RECT  2.350 0.865 2.470 1.270 ;
        END
        AntennaGateArea 0.088 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.435 -0.210 5.880 0.210 ;
        RECT  5.265 -0.210 5.435 0.595 ;
        RECT  4.685 -0.210 5.265 0.210 ;
        RECT  4.515 -0.210 4.685 0.715 ;
        RECT  2.270 -0.210 4.515 0.210 ;
        RECT  2.010 -0.210 2.270 0.300 ;
        RECT  1.430 -0.210 2.010 0.210 ;
        RECT  1.170 -0.210 1.430 0.415 ;
        RECT  0.265 -0.210 1.170 0.210 ;
        RECT  0.240 -0.210 0.265 0.285 ;
        RECT  0.120 -0.210 0.240 0.485 ;
        RECT  0.095 -0.210 0.120 0.285 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.425 2.310 5.880 2.730 ;
        RECT  5.165 2.015 5.425 2.730 ;
        RECT  4.440 2.310 5.165 2.730 ;
        RECT  4.270 2.055 4.440 2.730 ;
        RECT  3.400 2.310 4.270 2.730 ;
        RECT  3.140 2.020 3.400 2.730 ;
        RECT  2.610 2.310 3.140 2.730 ;
        RECT  2.350 1.965 2.610 2.730 ;
        RECT  1.285 2.310 2.350 2.730 ;
        RECT  1.165 1.995 1.285 2.730 ;
        RECT  0.265 2.310 1.165 2.730 ;
        RECT  0.095 1.650 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.880 2.520 ;
        LAYER M1 ;
        RECT  5.410 0.715 5.530 1.895 ;
        RECT  5.085 0.715 5.410 0.835 ;
        RECT  4.900 1.775 5.410 1.895 ;
        RECT  4.915 0.665 5.085 0.835 ;
        RECT  4.905 0.970 5.065 1.595 ;
        RECT  3.765 0.970 4.905 1.090 ;
        RECT  4.730 1.775 4.900 2.105 ;
        RECT  4.355 1.775 4.730 1.895 ;
        RECT  4.230 1.315 4.355 1.895 ;
        RECT  4.155 0.380 4.325 0.725 ;
        RECT  4.095 1.315 4.230 1.435 ;
        RECT  2.590 0.380 4.155 0.500 ;
        RECT  3.875 1.780 4.045 2.140 ;
        RECT  3.525 1.780 3.875 1.900 ;
        RECT  3.645 0.620 3.765 1.660 ;
        RECT  3.435 0.620 3.645 0.740 ;
        RECT  3.405 0.860 3.525 1.900 ;
        RECT  1.770 1.725 3.405 1.845 ;
        RECT  3.165 0.620 3.285 1.575 ;
        RECT  2.470 0.620 3.165 0.740 ;
        RECT  2.830 1.455 3.165 1.575 ;
        RECT  2.900 1.070 3.020 1.335 ;
        RECT  2.710 1.215 2.900 1.335 ;
        RECT  2.590 1.215 2.710 1.605 ;
        RECT  2.230 1.485 2.590 1.605 ;
        RECT  2.350 0.420 2.470 0.740 ;
        RECT  1.990 0.420 2.350 0.540 ;
        RECT  2.110 0.660 2.230 1.605 ;
        RECT  2.005 1.145 2.110 1.605 ;
        RECT  1.525 2.020 2.030 2.140 ;
        RECT  1.440 1.145 2.005 1.265 ;
        RECT  1.870 0.420 1.990 1.025 ;
        RECT  1.295 0.905 1.870 1.025 ;
        RECT  1.650 1.385 1.770 1.845 ;
        RECT  1.630 0.525 1.750 0.785 ;
        RECT  1.055 1.385 1.650 1.505 ;
        RECT  1.055 0.665 1.630 0.785 ;
        RECT  1.405 1.625 1.525 2.140 ;
        RECT  0.740 1.625 1.405 1.745 ;
        RECT  1.175 0.905 1.295 1.225 ;
        RECT  0.935 0.665 1.055 1.505 ;
        RECT  0.860 1.045 0.935 1.505 ;
        RECT  0.740 0.655 0.815 0.915 ;
        RECT  0.620 0.655 0.740 1.745 ;
    END
END DFFSQX2AD
MACRO DFFSQX4AD
    CLASS CORE ;
    FOREIGN DFFSQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.490 1.275 4.755 1.655 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.670 0.425 5.810 1.985 ;
        RECT  5.545 0.425 5.670 0.855 ;
        RECT  5.570 1.465 5.670 1.985 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.215 0.980 0.490 1.390 ;
        END
        AntennaGateArea 0.048 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.470 0.865 2.730 1.095 ;
        RECT  2.350 0.865 2.470 1.280 ;
        END
        AntennaGateArea 0.088 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.050 -0.210 6.160 0.210 ;
        RECT  5.930 -0.210 6.050 0.840 ;
        RECT  5.355 -0.210 5.930 0.210 ;
        RECT  5.185 -0.210 5.355 0.505 ;
        RECT  4.685 -0.210 5.185 0.210 ;
        RECT  4.515 -0.210 4.685 0.685 ;
        RECT  2.270 -0.210 4.515 0.210 ;
        RECT  2.010 -0.210 2.270 0.300 ;
        RECT  1.430 -0.210 2.010 0.210 ;
        RECT  1.170 -0.210 1.430 0.415 ;
        RECT  0.265 -0.210 1.170 0.210 ;
        RECT  0.095 -0.210 0.265 0.440 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.050 2.310 6.160 2.730 ;
        RECT  5.930 1.585 6.050 2.730 ;
        RECT  5.375 2.310 5.930 2.730 ;
        RECT  5.115 2.015 5.375 2.730 ;
        RECT  4.440 2.310 5.115 2.730 ;
        RECT  4.270 2.055 4.440 2.730 ;
        RECT  3.400 2.310 4.270 2.730 ;
        RECT  3.140 2.020 3.400 2.730 ;
        RECT  2.610 2.310 3.140 2.730 ;
        RECT  2.350 1.965 2.610 2.730 ;
        RECT  1.285 2.310 2.350 2.730 ;
        RECT  1.165 1.995 1.285 2.730 ;
        RECT  0.265 2.310 1.165 2.730 ;
        RECT  0.095 1.640 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.400 1.005 5.540 1.265 ;
        RECT  5.280 0.705 5.400 1.895 ;
        RECT  4.915 0.705 5.280 0.875 ;
        RECT  4.900 1.775 5.280 1.895 ;
        RECT  4.905 1.025 5.065 1.595 ;
        RECT  3.825 1.025 4.905 1.145 ;
        RECT  4.730 1.775 4.900 2.135 ;
        RECT  4.355 1.775 4.730 1.895 ;
        RECT  4.230 1.315 4.355 1.895 ;
        RECT  4.155 0.380 4.325 0.695 ;
        RECT  4.095 1.315 4.230 1.435 ;
        RECT  2.590 0.380 4.155 0.500 ;
        RECT  3.925 1.780 4.045 2.160 ;
        RECT  3.525 1.780 3.925 1.900 ;
        RECT  3.705 0.620 3.825 1.660 ;
        RECT  3.435 0.620 3.705 0.740 ;
        RECT  3.645 1.390 3.705 1.660 ;
        RECT  3.525 0.860 3.550 1.120 ;
        RECT  3.405 0.860 3.525 1.900 ;
        RECT  1.770 1.725 3.405 1.845 ;
        RECT  3.165 0.620 3.285 1.575 ;
        RECT  2.470 0.620 3.165 0.740 ;
        RECT  2.830 1.455 3.165 1.575 ;
        RECT  2.900 1.070 3.020 1.335 ;
        RECT  2.710 1.215 2.900 1.335 ;
        RECT  2.590 1.215 2.710 1.605 ;
        RECT  2.230 1.485 2.590 1.605 ;
        RECT  2.350 0.420 2.470 0.740 ;
        RECT  1.990 0.420 2.350 0.540 ;
        RECT  2.110 0.660 2.230 1.605 ;
        RECT  2.005 1.145 2.110 1.605 ;
        RECT  1.440 1.145 2.005 1.265 ;
        RECT  1.870 0.420 1.990 1.025 ;
        RECT  1.815 1.970 1.985 2.140 ;
        RECT  1.295 0.905 1.870 1.025 ;
        RECT  1.525 2.020 1.815 2.140 ;
        RECT  1.650 1.385 1.770 1.845 ;
        RECT  1.630 0.525 1.750 0.785 ;
        RECT  1.055 1.385 1.650 1.505 ;
        RECT  1.055 0.665 1.630 0.785 ;
        RECT  1.405 1.625 1.525 2.140 ;
        RECT  0.740 1.625 1.405 1.745 ;
        RECT  1.175 0.905 1.295 1.225 ;
        RECT  0.935 0.665 1.055 1.505 ;
        RECT  0.860 1.045 0.935 1.505 ;
        RECT  0.740 0.655 0.815 0.915 ;
        RECT  0.620 0.655 0.740 1.745 ;
    END
END DFFSQX4AD
MACRO DFFSQXLAD
    CLASS CORE ;
    FOREIGN DFFSQXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.475 1.305 4.735 1.685 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.410 0.360 5.530 1.685 ;
        RECT  5.335 0.360 5.410 0.530 ;
        RECT  5.370 1.425 5.410 1.685 ;
        END
        AntennaDiffArea 0.142 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 1.010 0.495 1.405 ;
        END
        AntennaGateArea 0.048 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.470 0.865 2.730 1.095 ;
        RECT  2.350 0.865 2.470 1.275 ;
        END
        AntennaGateArea 0.087 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.145 -0.210 5.600 0.210 ;
        RECT  4.975 -0.210 5.145 0.530 ;
        RECT  4.665 -0.210 4.975 0.210 ;
        RECT  4.495 -0.210 4.665 0.665 ;
        RECT  2.290 -0.210 4.495 0.210 ;
        RECT  2.030 -0.210 2.290 0.300 ;
        RECT  1.430 -0.210 2.030 0.210 ;
        RECT  1.170 -0.210 1.430 0.415 ;
        RECT  0.270 -0.210 1.170 0.210 ;
        RECT  0.100 -0.210 0.270 0.440 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.220 2.310 5.600 2.730 ;
        RECT  5.050 2.085 5.220 2.730 ;
        RECT  4.420 2.310 5.050 2.730 ;
        RECT  4.250 2.055 4.420 2.730 ;
        RECT  3.400 2.310 4.250 2.730 ;
        RECT  3.140 2.020 3.400 2.730 ;
        RECT  2.610 2.310 3.140 2.730 ;
        RECT  2.350 1.965 2.610 2.730 ;
        RECT  1.285 2.310 2.350 2.730 ;
        RECT  1.165 1.995 1.285 2.730 ;
        RECT  0.265 2.310 1.165 2.730 ;
        RECT  0.095 1.655 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  5.230 1.005 5.265 1.265 ;
        RECT  5.110 0.725 5.230 1.935 ;
        RECT  4.870 0.725 5.110 0.845 ;
        RECT  4.830 1.815 5.110 1.935 ;
        RECT  3.825 1.005 4.990 1.125 ;
        RECT  4.660 1.815 4.830 1.985 ;
        RECT  4.310 1.815 4.660 1.935 ;
        RECT  4.190 1.245 4.310 1.935 ;
        RECT  4.135 0.380 4.305 0.765 ;
        RECT  2.590 0.380 4.135 0.500 ;
        RECT  3.905 1.780 4.025 2.140 ;
        RECT  3.525 1.780 3.905 1.900 ;
        RECT  3.705 0.620 3.825 1.650 ;
        RECT  3.435 0.620 3.705 0.740 ;
        RECT  3.645 1.390 3.705 1.650 ;
        RECT  3.525 0.860 3.550 1.120 ;
        RECT  3.405 0.860 3.525 1.900 ;
        RECT  1.770 1.725 3.405 1.845 ;
        RECT  3.165 0.620 3.285 1.575 ;
        RECT  2.470 0.620 3.165 0.740 ;
        RECT  2.830 1.455 3.165 1.575 ;
        RECT  2.900 1.070 3.020 1.335 ;
        RECT  2.710 1.215 2.900 1.335 ;
        RECT  2.590 1.215 2.710 1.605 ;
        RECT  2.230 1.485 2.590 1.605 ;
        RECT  2.350 0.420 2.470 0.740 ;
        RECT  1.990 0.420 2.350 0.540 ;
        RECT  2.110 0.660 2.230 1.605 ;
        RECT  2.005 1.145 2.110 1.605 ;
        RECT  1.525 1.970 2.030 2.140 ;
        RECT  1.440 1.145 2.005 1.265 ;
        RECT  1.870 0.420 1.990 1.025 ;
        RECT  1.295 0.905 1.870 1.025 ;
        RECT  1.650 1.385 1.770 1.845 ;
        RECT  1.630 0.525 1.750 0.785 ;
        RECT  1.055 1.385 1.650 1.505 ;
        RECT  1.055 0.665 1.630 0.785 ;
        RECT  1.405 1.625 1.525 2.140 ;
        RECT  0.740 1.625 1.405 1.745 ;
        RECT  1.175 0.905 1.295 1.225 ;
        RECT  0.935 0.665 1.055 1.505 ;
        RECT  0.860 1.045 0.935 1.505 ;
        RECT  0.740 0.655 0.815 0.915 ;
        RECT  0.620 0.655 0.740 1.745 ;
    END
END DFFSQXLAD
MACRO DFFSRHQX1AD
    CLASS CORE ;
    FOREIGN DFFSRHQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.585 1.050 2.860 1.375 ;
        RECT  2.540 1.080 2.585 1.200 ;
        END
        AntennaGateArea 0.111 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.975 1.020 7.095 1.280 ;
        RECT  5.810 1.080 6.975 1.200 ;
        RECT  5.670 1.080 5.810 1.375 ;
        END
        AntennaGateArea 0.101 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.130 1.145 9.170 1.375 ;
        RECT  9.010 0.645 9.130 1.935 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.710 0.985 1.925 1.375 ;
        END
        AntennaGateArea 0.05 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.930 0.495 1.375 ;
        END
        AntennaGateArea 0.12 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.800 -0.210 9.240 0.210 ;
        RECT  8.540 -0.210 8.800 0.310 ;
        RECT  7.595 -0.210 8.540 0.210 ;
        RECT  7.335 -0.210 7.595 0.310 ;
        RECT  5.835 -0.210 7.335 0.210 ;
        RECT  5.575 -0.210 5.835 0.300 ;
        RECT  4.605 -0.210 5.575 0.210 ;
        RECT  4.345 -0.210 4.605 0.300 ;
        RECT  2.745 -0.210 4.345 0.210 ;
        RECT  2.485 -0.210 2.745 0.300 ;
        RECT  1.755 -0.210 2.485 0.210 ;
        RECT  1.495 -0.210 1.755 0.300 ;
        RECT  0.680 -0.210 1.495 0.210 ;
        RECT  0.420 -0.210 0.680 0.300 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.810 2.310 9.240 2.730 ;
        RECT  8.550 2.005 8.810 2.730 ;
        RECT  7.445 2.310 8.550 2.730 ;
        RECT  7.185 2.220 7.445 2.730 ;
        RECT  5.755 2.310 7.185 2.730 ;
        RECT  5.495 2.225 5.755 2.730 ;
        RECT  5.005 2.310 5.495 2.730 ;
        RECT  4.745 2.225 5.005 2.730 ;
        RECT  4.215 2.310 4.745 2.730 ;
        RECT  3.955 2.225 4.215 2.730 ;
        RECT  2.775 2.310 3.955 2.730 ;
        RECT  2.515 2.225 2.775 2.730 ;
        RECT  1.895 2.310 2.515 2.730 ;
        RECT  1.635 2.225 1.895 2.730 ;
        RECT  0.575 2.310 1.635 2.730 ;
        RECT  0.355 1.880 0.575 2.730 ;
        RECT  0.000 2.310 0.355 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.240 2.520 ;
        LAYER M1 ;
        RECT  8.775 1.000 8.880 1.260 ;
        RECT  8.655 0.430 8.775 1.885 ;
        RECT  6.705 0.430 8.655 0.550 ;
        RECT  8.500 1.000 8.655 1.260 ;
        RECT  8.285 1.765 8.655 1.885 ;
        RECT  8.380 0.695 8.410 0.905 ;
        RECT  8.215 0.695 8.380 1.590 ;
        RECT  8.025 1.765 8.285 2.045 ;
        RECT  7.575 0.695 8.215 0.815 ;
        RECT  7.955 1.160 8.075 1.645 ;
        RECT  6.535 1.925 8.025 2.045 ;
        RECT  7.335 1.160 7.955 1.280 ;
        RECT  6.920 1.400 7.835 1.575 ;
        RECT  7.455 0.695 7.575 1.040 ;
        RECT  7.215 0.780 7.335 1.280 ;
        RECT  6.325 0.780 7.215 0.900 ;
        RECT  6.705 1.400 6.920 1.805 ;
        RECT  6.445 0.430 6.705 0.660 ;
        RECT  6.320 1.675 6.705 1.805 ;
        RECT  6.050 1.435 6.415 1.555 ;
        RECT  6.205 0.420 6.325 0.900 ;
        RECT  6.170 1.675 6.320 1.865 ;
        RECT  5.965 1.985 6.225 2.165 ;
        RECT  3.955 0.420 6.205 0.540 ;
        RECT  4.795 1.745 6.170 1.865 ;
        RECT  5.070 0.680 6.085 0.805 ;
        RECT  5.930 1.435 6.050 1.615 ;
        RECT  4.585 1.985 5.965 2.105 ;
        RECT  5.070 1.495 5.930 1.615 ;
        RECT  4.915 0.680 5.070 1.615 ;
        RECT  4.675 0.660 4.795 1.865 ;
        RECT  2.415 0.660 4.675 0.780 ;
        RECT  4.325 1.985 4.585 2.170 ;
        RECT  4.420 0.900 4.495 1.160 ;
        RECT  4.250 0.900 4.420 1.835 ;
        RECT  3.275 1.985 4.325 2.105 ;
        RECT  3.465 0.900 4.250 1.080 ;
        RECT  3.515 1.715 4.250 1.835 ;
        RECT  3.695 0.380 3.955 0.540 ;
        RECT  1.785 0.420 3.695 0.540 ;
        RECT  3.395 1.540 3.515 1.835 ;
        RECT  3.155 0.990 3.275 2.105 ;
        RECT  3.065 0.990 3.155 1.250 ;
        RECT  1.155 1.985 3.155 2.105 ;
        RECT  2.175 1.740 3.035 1.860 ;
        RECT  2.295 0.660 2.415 1.590 ;
        RECT  2.045 0.660 2.175 1.860 ;
        RECT  1.920 0.660 2.045 0.830 ;
        RECT  1.915 1.740 2.045 1.860 ;
        RECT  1.665 0.420 1.785 0.815 ;
        RECT  1.260 0.695 1.665 0.815 ;
        RECT  1.260 1.390 1.505 1.510 ;
        RECT  1.205 0.330 1.375 0.540 ;
        RECT  1.115 0.695 1.260 1.510 ;
        RECT  0.230 0.420 1.205 0.540 ;
        RECT  0.990 1.670 1.155 2.105 ;
        RECT  0.890 1.095 1.115 1.270 ;
        RECT  0.870 1.460 0.990 2.105 ;
        RECT  0.770 0.660 0.905 0.920 ;
        RECT  0.770 1.460 0.870 1.580 ;
        RECT  0.650 0.660 0.770 1.580 ;
        RECT  0.110 0.420 0.230 1.610 ;
    END
END DFFSRHQX1AD
MACRO DFFSRHQX2AD
    CLASS CORE ;
    FOREIGN DFFSRHQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.585 1.050 2.860 1.375 ;
        RECT  2.540 1.080 2.585 1.200 ;
        END
        AntennaGateArea 0.131 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.975 1.020 7.095 1.280 ;
        RECT  5.810 1.080 6.975 1.200 ;
        RECT  5.670 1.080 5.810 1.375 ;
        END
        AntennaGateArea 0.131 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.130 1.145 9.170 1.375 ;
        RECT  9.010 0.370 9.130 1.990 ;
        END
        AntennaDiffArea 0.365 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.710 0.985 1.925 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.930 0.495 1.375 ;
        END
        AntennaGateArea 0.116 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.770 -0.210 9.240 0.210 ;
        RECT  8.510 -0.210 8.770 0.310 ;
        RECT  7.595 -0.210 8.510 0.210 ;
        RECT  7.335 -0.210 7.595 0.310 ;
        RECT  5.835 -0.210 7.335 0.210 ;
        RECT  5.575 -0.210 5.835 0.300 ;
        RECT  4.605 -0.210 5.575 0.210 ;
        RECT  4.345 -0.210 4.605 0.300 ;
        RECT  2.745 -0.210 4.345 0.210 ;
        RECT  2.485 -0.210 2.745 0.300 ;
        RECT  1.755 -0.210 2.485 0.210 ;
        RECT  1.495 -0.210 1.755 0.300 ;
        RECT  0.680 -0.210 1.495 0.210 ;
        RECT  0.420 -0.210 0.680 0.300 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.810 2.310 9.240 2.730 ;
        RECT  8.550 2.010 8.810 2.730 ;
        RECT  7.445 2.310 8.550 2.730 ;
        RECT  7.185 2.220 7.445 2.730 ;
        RECT  5.755 2.310 7.185 2.730 ;
        RECT  5.495 2.230 5.755 2.730 ;
        RECT  5.005 2.310 5.495 2.730 ;
        RECT  4.745 2.230 5.005 2.730 ;
        RECT  4.215 2.310 4.745 2.730 ;
        RECT  3.955 2.230 4.215 2.730 ;
        RECT  2.775 2.310 3.955 2.730 ;
        RECT  2.515 2.230 2.775 2.730 ;
        RECT  1.895 2.310 2.515 2.730 ;
        RECT  1.635 2.230 1.895 2.730 ;
        RECT  0.575 2.310 1.635 2.730 ;
        RECT  0.355 1.880 0.575 2.730 ;
        RECT  0.000 2.310 0.355 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.240 2.520 ;
        LAYER M1 ;
        RECT  8.775 1.000 8.880 1.260 ;
        RECT  8.655 0.430 8.775 1.885 ;
        RECT  6.705 0.430 8.655 0.550 ;
        RECT  8.500 1.000 8.655 1.260 ;
        RECT  8.285 1.765 8.655 1.885 ;
        RECT  8.380 0.695 8.410 0.905 ;
        RECT  8.215 0.695 8.380 1.590 ;
        RECT  8.025 1.765 8.285 2.045 ;
        RECT  7.575 0.695 8.215 0.815 ;
        RECT  7.955 1.160 8.075 1.645 ;
        RECT  6.535 1.925 8.025 2.045 ;
        RECT  7.335 1.160 7.955 1.280 ;
        RECT  6.895 1.400 7.835 1.575 ;
        RECT  7.455 0.695 7.575 1.040 ;
        RECT  7.215 0.780 7.335 1.280 ;
        RECT  6.325 0.780 7.215 0.900 ;
        RECT  6.705 1.400 6.895 1.805 ;
        RECT  6.445 0.430 6.705 0.660 ;
        RECT  6.320 1.675 6.705 1.805 ;
        RECT  6.050 1.435 6.415 1.555 ;
        RECT  6.205 0.420 6.325 0.900 ;
        RECT  6.170 1.675 6.320 1.865 ;
        RECT  5.965 1.990 6.225 2.190 ;
        RECT  3.955 0.420 6.205 0.540 ;
        RECT  4.795 1.745 6.170 1.865 ;
        RECT  5.070 0.680 6.085 0.805 ;
        RECT  5.930 1.435 6.050 1.615 ;
        RECT  4.585 1.990 5.965 2.110 ;
        RECT  5.070 1.495 5.930 1.615 ;
        RECT  4.915 0.680 5.070 1.615 ;
        RECT  4.675 0.660 4.795 1.865 ;
        RECT  2.415 0.660 4.675 0.780 ;
        RECT  4.325 1.990 4.585 2.170 ;
        RECT  4.420 0.900 4.495 1.160 ;
        RECT  4.420 1.690 4.465 1.810 ;
        RECT  4.250 0.900 4.420 1.835 ;
        RECT  3.275 1.990 4.325 2.110 ;
        RECT  3.465 0.900 4.250 1.080 ;
        RECT  4.205 1.690 4.250 1.835 ;
        RECT  3.515 1.715 4.205 1.835 ;
        RECT  3.695 0.380 3.955 0.540 ;
        RECT  1.785 0.420 3.695 0.540 ;
        RECT  3.395 1.540 3.515 1.835 ;
        RECT  3.155 0.990 3.275 2.110 ;
        RECT  3.065 0.990 3.155 1.250 ;
        RECT  1.155 1.990 3.155 2.110 ;
        RECT  2.175 1.740 3.035 1.860 ;
        RECT  2.295 0.660 2.415 1.590 ;
        RECT  2.045 0.670 2.175 1.860 ;
        RECT  1.920 0.670 2.045 0.840 ;
        RECT  1.915 1.740 2.045 1.860 ;
        RECT  1.665 0.420 1.785 0.815 ;
        RECT  1.260 0.695 1.665 0.815 ;
        RECT  1.260 1.390 1.505 1.510 ;
        RECT  1.115 0.335 1.375 0.540 ;
        RECT  1.115 0.695 1.260 1.510 ;
        RECT  0.990 1.675 1.155 2.110 ;
        RECT  0.230 0.420 1.115 0.540 ;
        RECT  0.890 1.095 1.115 1.270 ;
        RECT  0.870 1.460 0.990 2.110 ;
        RECT  0.770 0.660 0.905 0.920 ;
        RECT  0.770 1.460 0.870 1.580 ;
        RECT  0.650 0.660 0.770 1.580 ;
        RECT  0.110 0.420 0.230 1.610 ;
    END
END DFFSRHQX2AD
MACRO DFFSRHQX4AD
    CLASS CORE ;
    FOREIGN DFFSRHQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.865 1.050 3.140 1.375 ;
        RECT  2.820 1.080 2.865 1.200 ;
        END
        AntennaGateArea 0.159 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.310 1.025 9.455 1.330 ;
        RECT  8.090 1.190 9.310 1.330 ;
        RECT  7.925 1.190 8.090 1.380 ;
        RECT  7.240 1.260 7.925 1.380 ;
        END
        AntennaGateArea 0.215 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.270 0.355 11.410 2.040 ;
        RECT  11.170 0.355 11.270 0.875 ;
        RECT  11.170 1.520 11.270 2.040 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 0.865 2.215 1.125 ;
        END
        AntennaGateArea 0.072 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.930 0.490 1.375 ;
        END
        AntennaGateArea 0.172 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.650 -0.210 11.760 0.210 ;
        RECT  11.530 -0.210 11.650 0.875 ;
        RECT  10.845 -0.210 11.530 0.210 ;
        RECT  10.585 -0.210 10.845 0.310 ;
        RECT  9.900 -0.210 10.585 0.210 ;
        RECT  9.730 -0.210 9.900 0.260 ;
        RECT  7.145 -0.210 9.730 0.210 ;
        RECT  6.885 -0.210 7.145 0.630 ;
        RECT  5.935 -0.210 6.885 0.210 ;
        RECT  5.675 -0.210 5.935 0.300 ;
        RECT  4.995 -0.210 5.675 0.210 ;
        RECT  4.735 -0.210 4.995 0.300 ;
        RECT  3.010 -0.210 4.735 0.210 ;
        RECT  2.840 -0.210 3.010 0.260 ;
        RECT  2.000 -0.210 2.840 0.210 ;
        RECT  1.830 -0.210 2.000 0.260 ;
        RECT  0.545 -0.210 1.830 0.210 ;
        RECT  0.375 -0.210 0.545 0.260 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.650 2.310 11.760 2.730 ;
        RECT  11.530 1.590 11.650 2.730 ;
        RECT  10.980 2.310 11.530 2.730 ;
        RECT  10.720 2.010 10.980 2.730 ;
        RECT  9.560 2.310 10.720 2.730 ;
        RECT  9.300 2.210 9.560 2.730 ;
        RECT  6.905 2.310 9.300 2.730 ;
        RECT  6.475 2.260 6.905 2.730 ;
        RECT  5.825 2.310 6.475 2.730 ;
        RECT  5.655 2.260 5.825 2.730 ;
        RECT  4.565 2.310 5.655 2.730 ;
        RECT  4.305 1.890 4.565 2.730 ;
        RECT  3.055 2.310 4.305 2.730 ;
        RECT  2.795 2.220 3.055 2.730 ;
        RECT  2.140 2.310 2.795 2.730 ;
        RECT  1.970 2.265 2.140 2.730 ;
        RECT  1.380 2.310 1.970 2.730 ;
        RECT  1.210 2.265 1.380 2.730 ;
        RECT  0.570 2.310 1.210 2.730 ;
        RECT  0.350 2.050 0.570 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.760 2.520 ;
        LAYER M1 ;
        RECT  10.940 1.000 11.105 1.260 ;
        RECT  10.820 0.470 10.940 1.890 ;
        RECT  10.240 0.470 10.820 0.590 ;
        RECT  10.725 1.000 10.820 1.260 ;
        RECT  10.480 1.770 10.820 1.890 ;
        RECT  10.605 0.710 10.630 0.905 ;
        RECT  10.485 0.710 10.605 1.590 ;
        RECT  10.460 0.710 10.485 0.905 ;
        RECT  10.310 1.770 10.480 2.085 ;
        RECT  9.935 0.710 10.460 0.835 ;
        RECT  10.160 1.090 10.330 1.635 ;
        RECT  9.150 1.965 10.310 2.085 ;
        RECT  10.070 0.350 10.240 0.590 ;
        RECT  9.695 1.090 10.160 1.210 ;
        RECT  8.045 0.380 10.070 0.500 ;
        RECT  9.885 1.360 10.005 1.620 ;
        RECT  9.815 0.710 9.935 0.970 ;
        RECT  8.910 1.460 9.885 1.580 ;
        RECT  9.575 0.660 9.695 1.210 ;
        RECT  7.455 0.660 9.575 0.780 ;
        RECT  9.030 1.965 9.150 2.140 ;
        RECT  8.000 2.020 9.030 2.140 ;
        RECT  8.790 1.460 8.910 1.900 ;
        RECT  7.130 1.780 8.790 1.900 ;
        RECT  7.825 0.900 8.685 1.020 ;
        RECT  7.730 1.540 8.650 1.660 ;
        RECT  7.625 0.900 7.825 1.110 ;
        RECT  7.470 1.500 7.730 1.660 ;
        RECT  5.455 2.020 7.710 2.140 ;
        RECT  6.465 0.990 7.625 1.110 ;
        RECT  6.465 1.500 7.470 1.620 ;
        RECT  7.335 0.660 7.455 0.870 ;
        RECT  6.705 0.750 7.335 0.870 ;
        RECT  7.010 1.740 7.130 1.900 ;
        RECT  5.420 1.740 7.010 1.860 ;
        RECT  6.585 0.420 6.705 0.870 ;
        RECT  5.385 0.420 6.585 0.540 ;
        RECT  6.345 0.660 6.465 1.620 ;
        RECT  6.010 1.385 6.345 1.620 ;
        RECT  6.085 0.660 6.205 1.260 ;
        RECT  2.695 0.660 6.085 0.780 ;
        RECT  5.420 1.140 6.085 1.260 ;
        RECT  5.540 1.385 6.010 1.505 ;
        RECT  5.075 0.900 5.965 1.020 ;
        RECT  5.195 2.020 5.455 2.185 ;
        RECT  5.300 1.140 5.420 1.860 ;
        RECT  5.125 0.340 5.385 0.540 ;
        RECT  4.805 2.020 5.195 2.140 ;
        RECT  5.075 1.635 5.180 1.895 ;
        RECT  3.100 0.420 5.125 0.540 ;
        RECT  4.955 0.900 5.075 1.895 ;
        RECT  3.735 0.900 4.955 1.020 ;
        RECT  3.795 1.405 4.955 1.525 ;
        RECT  4.685 1.645 4.805 2.140 ;
        RECT  4.035 1.645 4.685 1.765 ;
        RECT  3.555 1.140 4.510 1.260 ;
        RECT  3.915 1.645 4.035 2.125 ;
        RECT  3.555 2.005 3.915 2.125 ;
        RECT  3.675 1.405 3.795 1.885 ;
        RECT  3.435 0.990 3.555 2.125 ;
        RECT  3.345 0.990 3.435 1.260 ;
        RECT  1.240 1.980 3.435 2.100 ;
        RECT  2.455 1.740 3.315 1.860 ;
        RECT  2.980 0.380 3.100 0.540 ;
        RECT  1.805 0.380 2.980 0.500 ;
        RECT  2.575 0.660 2.695 1.590 ;
        RECT  2.335 0.620 2.455 1.860 ;
        RECT  2.165 0.620 2.335 0.740 ;
        RECT  2.235 1.740 2.335 1.860 ;
        RECT  1.685 0.380 1.805 1.740 ;
        RECT  1.450 0.595 1.685 0.780 ;
        RECT  1.545 1.620 1.685 1.740 ;
        RECT  1.260 0.660 1.450 0.780 ;
        RECT  1.330 0.330 1.405 0.450 ;
        RECT  1.145 0.330 1.330 0.500 ;
        RECT  1.090 0.660 1.260 1.090 ;
        RECT  0.980 1.260 1.240 2.100 ;
        RECT  0.230 0.380 1.145 0.500 ;
        RECT  0.730 1.260 0.980 1.380 ;
        RECT  0.730 0.620 0.970 0.740 ;
        RECT  0.610 0.620 0.730 1.380 ;
        RECT  0.110 0.380 0.230 1.600 ;
    END
END DFFSRHQX4AD
MACRO DFFSRHQX8AD
    CLASS CORE ;
    FOREIGN DFFSRHQX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.070 1.070 3.305 1.375 ;
        END
        AntennaGateArea 0.233 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.715 0.925 9.835 1.220 ;
        RECT  8.235 1.100 9.715 1.220 ;
        RECT  7.725 1.100 8.235 1.330 ;
        RECT  7.110 1.100 7.725 1.220 ;
        RECT  6.940 0.965 7.110 1.220 ;
        END
        AntennaGateArea 0.272 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.545 0.365 12.715 2.165 ;
        RECT  11.995 1.050 12.545 1.475 ;
        RECT  11.785 0.365 11.995 2.165 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.980 2.315 1.375 ;
        END
        AntennaGateArea 0.139 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.025 0.550 1.405 ;
        END
        AntennaGateArea 0.265 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.075 -0.210 13.160 0.210 ;
        RECT  12.905 -0.210 13.075 0.795 ;
        RECT  12.355 -0.210 12.905 0.210 ;
        RECT  12.185 -0.210 12.355 0.795 ;
        RECT  11.610 -0.210 12.185 0.210 ;
        RECT  11.350 -0.210 11.610 0.310 ;
        RECT  10.445 -0.210 11.350 0.210 ;
        RECT  10.185 -0.210 10.445 0.310 ;
        RECT  8.185 -0.210 10.185 0.210 ;
        RECT  8.065 -0.210 8.185 0.500 ;
        RECT  7.015 -0.210 8.065 0.210 ;
        RECT  6.755 -0.210 7.015 0.260 ;
        RECT  6.265 -0.210 6.755 0.210 ;
        RECT  5.745 -0.210 6.265 0.260 ;
        RECT  3.250 -0.210 5.745 0.210 ;
        RECT  2.990 -0.210 3.250 0.310 ;
        RECT  1.990 -0.210 2.990 0.210 ;
        RECT  1.730 -0.210 1.990 0.310 ;
        RECT  0.680 -0.210 1.730 0.210 ;
        RECT  0.420 -0.210 0.680 0.250 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.075 2.310 13.160 2.730 ;
        RECT  12.905 1.475 13.075 2.730 ;
        RECT  12.355 2.310 12.905 2.730 ;
        RECT  12.185 1.735 12.355 2.730 ;
        RECT  11.610 2.310 12.185 2.730 ;
        RECT  11.350 2.220 11.610 2.730 ;
        RECT  10.170 2.310 11.350 2.730 ;
        RECT  9.910 2.220 10.170 2.730 ;
        RECT  7.495 2.310 9.910 2.730 ;
        RECT  7.235 2.260 7.495 2.730 ;
        RECT  6.565 2.310 7.235 2.730 ;
        RECT  6.305 2.260 6.565 2.730 ;
        RECT  5.095 2.310 6.305 2.730 ;
        RECT  4.835 2.260 5.095 2.730 ;
        RECT  3.415 2.310 4.835 2.730 ;
        RECT  3.155 2.290 3.415 2.730 ;
        RECT  2.295 2.310 3.155 2.730 ;
        RECT  2.035 2.260 2.295 2.730 ;
        RECT  1.490 2.310 2.035 2.730 ;
        RECT  1.320 2.185 1.490 2.730 ;
        RECT  0.540 2.310 1.320 2.730 ;
        RECT  0.370 2.245 0.540 2.730 ;
        RECT  0.000 2.310 0.370 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 13.160 2.520 ;
        LAYER M1 ;
        RECT  11.545 1.060 11.665 1.230 ;
        RECT  11.395 0.430 11.545 2.100 ;
        RECT  9.795 0.430 11.395 0.550 ;
        RECT  11.235 1.060 11.395 1.230 ;
        RECT  11.055 1.970 11.395 2.100 ;
        RECT  11.100 0.670 11.160 0.950 ;
        RECT  11.100 1.375 11.105 1.545 ;
        RECT  10.980 0.670 11.100 1.545 ;
        RECT  10.795 1.780 11.055 2.100 ;
        RECT  10.315 0.670 10.980 0.790 ;
        RECT  10.935 1.375 10.980 1.545 ;
        RECT  10.695 1.130 10.815 1.660 ;
        RECT  8.380 1.980 10.795 2.100 ;
        RECT  10.075 1.130 10.695 1.250 ;
        RECT  10.375 1.400 10.495 1.660 ;
        RECT  9.365 1.400 10.375 1.520 ;
        RECT  10.195 0.670 10.315 1.000 ;
        RECT  9.955 0.670 10.075 1.250 ;
        RECT  9.585 0.670 9.955 0.790 ;
        RECT  9.690 0.380 9.795 0.550 ;
        RECT  8.445 0.380 9.690 0.500 ;
        RECT  9.455 0.620 9.585 0.790 ;
        RECT  7.885 0.620 9.455 0.740 ;
        RECT  9.245 1.400 9.365 1.860 ;
        RECT  7.930 1.740 9.245 1.860 ;
        RECT  7.645 0.860 9.095 0.980 ;
        RECT  7.285 1.500 9.000 1.620 ;
        RECT  7.825 2.015 8.085 2.190 ;
        RECT  7.810 1.740 7.930 1.895 ;
        RECT  7.765 0.380 7.885 0.740 ;
        RECT  5.965 2.015 7.825 2.140 ;
        RECT  6.050 1.775 7.810 1.895 ;
        RECT  5.580 0.380 7.765 0.500 ;
        RECT  7.525 0.620 7.645 0.980 ;
        RECT  6.685 0.620 7.525 0.740 ;
        RECT  7.165 1.500 7.285 1.655 ;
        RECT  6.685 1.535 7.165 1.655 ;
        RECT  6.565 0.620 6.685 1.655 ;
        RECT  6.170 1.410 6.565 1.530 ;
        RECT  6.305 0.620 6.425 1.285 ;
        RECT  3.725 0.620 6.305 0.740 ;
        RECT  6.050 1.165 6.305 1.285 ;
        RECT  5.810 0.925 6.165 1.045 ;
        RECT  5.930 1.165 6.050 1.895 ;
        RECT  5.705 2.015 5.965 2.190 ;
        RECT  5.690 0.925 5.810 1.850 ;
        RECT  3.945 2.015 5.705 2.140 ;
        RECT  5.100 0.925 5.690 1.045 ;
        RECT  4.125 1.730 5.690 1.850 ;
        RECT  5.320 0.335 5.580 0.500 ;
        RECT  5.405 1.325 5.525 1.585 ;
        RECT  4.265 1.410 5.405 1.530 ;
        RECT  3.480 0.380 5.320 0.500 ;
        RECT  4.980 0.870 5.100 1.045 ;
        RECT  4.005 0.870 4.980 0.990 ;
        RECT  3.945 1.110 4.775 1.230 ;
        RECT  3.855 1.110 3.945 2.140 ;
        RECT  3.825 1.090 3.855 2.140 ;
        RECT  3.495 1.090 3.825 1.230 ;
        RECT  2.215 2.020 3.825 2.140 ;
        RECT  3.590 0.620 3.725 0.795 ;
        RECT  2.630 1.780 3.680 1.900 ;
        RECT  2.950 0.675 3.590 0.795 ;
        RECT  3.360 0.380 3.480 0.550 ;
        RECT  1.895 0.430 3.360 0.550 ;
        RECT  2.950 1.540 3.015 1.660 ;
        RECT  2.830 0.675 2.950 1.660 ;
        RECT  2.680 0.675 2.830 0.935 ;
        RECT  2.755 1.540 2.830 1.660 ;
        RECT  2.560 1.425 2.630 1.900 ;
        RECT  2.440 0.670 2.560 1.900 ;
        RECT  2.260 0.670 2.440 0.790 ;
        RECT  2.095 1.925 2.215 2.140 ;
        RECT  1.220 1.925 2.095 2.045 ;
        RECT  1.775 0.430 1.895 0.855 ;
        RECT  1.725 1.160 1.845 1.715 ;
        RECT  1.475 0.735 1.775 0.855 ;
        RECT  1.475 1.160 1.725 1.280 ;
        RECT  1.305 0.735 1.475 1.280 ;
        RECT  0.240 0.380 1.320 0.500 ;
        RECT  0.980 1.160 1.305 1.280 ;
        RECT  1.050 1.575 1.220 2.045 ;
        RECT  0.790 1.575 1.050 1.695 ;
        RECT  0.870 0.690 0.990 0.950 ;
        RECT  0.790 0.830 0.870 0.950 ;
        RECT  0.670 0.830 0.790 1.695 ;
        RECT  0.205 1.555 0.255 1.985 ;
        RECT  0.205 0.380 0.240 0.900 ;
        RECT  0.085 0.380 0.205 1.985 ;
    END
END DFFSRHQX8AD
MACRO DFFSRX1AD
    CLASS CORE ;
    FOREIGN DFFSRX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.185 0.960 6.420 1.395 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.980 3.010 1.440 ;
        END
        AntennaGateArea 0.048 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.290 1.360 7.490 1.655 ;
        RECT  7.125 0.680 7.290 1.655 ;
        END
        AntennaDiffArea 0.207 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.890 0.615 8.050 1.890 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.180 1.050 0.490 1.420 ;
        END
        AntennaGateArea 0.048 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.585 1.025 2.730 1.540 ;
        END
        AntennaGateArea 0.083 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.675 -0.210 8.120 0.210 ;
        RECT  7.505 -0.210 7.675 0.825 ;
        RECT  6.605 -0.210 7.505 0.210 ;
        RECT  6.435 -0.210 6.605 0.525 ;
        RECT  2.850 -0.210 6.435 0.210 ;
        RECT  2.590 -0.210 2.850 0.300 ;
        RECT  1.620 -0.210 2.590 0.210 ;
        RECT  1.450 -0.210 1.620 0.605 ;
        RECT  0.340 -0.210 1.450 0.210 ;
        RECT  0.170 -0.210 0.340 0.850 ;
        RECT  0.000 -0.210 0.170 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.700 2.310 8.120 2.730 ;
        RECT  7.440 2.015 7.700 2.730 ;
        RECT  6.965 2.310 7.440 2.730 ;
        RECT  6.705 2.015 6.965 2.730 ;
        RECT  5.020 2.310 6.705 2.730 ;
        RECT  4.760 2.210 5.020 2.730 ;
        RECT  3.480 2.310 4.760 2.730 ;
        RECT  3.220 2.040 3.480 2.730 ;
        RECT  2.820 2.310 3.220 2.730 ;
        RECT  2.560 2.075 2.820 2.730 ;
        RECT  1.560 2.310 2.560 2.730 ;
        RECT  1.440 1.995 1.560 2.730 ;
        RECT  0.340 2.310 1.440 2.730 ;
        RECT  0.170 1.685 0.340 2.730 ;
        RECT  0.000 2.310 0.170 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.120 2.520 ;
        LAYER M1 ;
        RECT  7.650 1.020 7.770 1.895 ;
        RECT  7.005 1.775 7.650 1.895 ;
        RECT  6.885 0.355 7.005 1.895 ;
        RECT  6.795 0.355 6.885 0.525 ;
        RECT  5.790 1.535 6.885 1.710 ;
        RECT  6.605 0.670 6.725 1.365 ;
        RECT  4.870 0.670 6.605 0.790 ;
        RECT  4.115 0.380 6.290 0.500 ;
        RECT  5.870 1.855 6.130 2.090 ;
        RECT  3.620 1.970 5.870 2.090 ;
        RECT  5.435 0.960 5.605 1.850 ;
        RECT  5.185 0.960 5.435 1.115 ;
        RECT  3.490 1.730 5.435 1.850 ;
        RECT  4.870 1.480 5.295 1.600 ;
        RECT  4.750 0.670 4.870 1.600 ;
        RECT  4.510 0.830 4.630 1.600 ;
        RECT  4.370 0.830 4.510 1.010 ;
        RECT  4.060 1.480 4.510 1.600 ;
        RECT  3.635 1.200 4.385 1.320 ;
        RECT  3.875 0.890 4.370 1.010 ;
        RECT  3.995 0.380 4.115 0.770 ;
        RECT  3.755 0.420 3.875 1.010 ;
        RECT  2.225 0.420 3.755 0.540 ;
        RECT  3.515 0.660 3.635 1.320 ;
        RECT  2.490 0.660 3.515 0.780 ;
        RECT  3.370 1.730 3.490 1.920 ;
        RECT  3.315 0.900 3.390 1.020 ;
        RECT  2.845 1.800 3.370 1.920 ;
        RECT  3.250 0.900 3.315 1.430 ;
        RECT  3.130 0.900 3.250 1.680 ;
        RECT  2.970 1.560 3.130 1.680 ;
        RECT  2.725 1.730 2.845 1.920 ;
        RECT  2.040 1.730 2.725 1.850 ;
        RECT  2.465 0.660 2.490 0.920 ;
        RECT  2.345 0.660 2.465 1.610 ;
        RECT  2.175 1.255 2.345 1.610 ;
        RECT  2.105 0.420 2.225 1.135 ;
        RECT  1.800 2.020 2.200 2.140 ;
        RECT  1.595 1.255 2.175 1.375 ;
        RECT  1.405 1.015 2.105 1.135 ;
        RECT  1.920 1.515 2.040 1.850 ;
        RECT  1.865 0.635 1.985 0.895 ;
        RECT  1.165 1.515 1.920 1.635 ;
        RECT  1.165 0.775 1.865 0.895 ;
        RECT  1.680 1.755 1.800 2.140 ;
        RECT  0.835 1.755 1.680 1.875 ;
        RECT  1.285 1.015 1.405 1.285 ;
        RECT  1.045 0.775 1.165 1.635 ;
        RECT  0.955 1.175 1.045 1.635 ;
        RECT  0.835 0.635 0.925 0.895 ;
        RECT  0.715 0.635 0.835 1.875 ;
    END
END DFFSRX1AD
MACRO DFFSRX2AD
    CLASS CORE ;
    FOREIGN DFFSRX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.465 0.955 6.700 1.395 ;
        END
        AntennaGateArea 0.101 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.880 3.010 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.570 1.360 7.770 1.655 ;
        RECT  7.405 0.415 7.570 1.655 ;
        END
        AntennaDiffArea 0.373 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.290 0.615 8.330 1.985 ;
        RECT  8.170 0.415 8.290 1.985 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 1.375 0.535 1.700 ;
        END
        AntennaGateArea 0.048 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.565 0.990 2.730 1.540 ;
        END
        AntennaGateArea 0.096 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.955 -0.210 8.400 0.210 ;
        RECT  7.785 -0.210 7.955 0.810 ;
        RECT  6.885 -0.210 7.785 0.210 ;
        RECT  6.715 -0.210 6.885 0.525 ;
        RECT  2.885 -0.210 6.715 0.210 ;
        RECT  2.625 -0.210 2.885 0.260 ;
        RECT  1.585 -0.210 2.625 0.210 ;
        RECT  1.415 -0.210 1.585 0.650 ;
        RECT  0.295 -0.210 1.415 0.210 ;
        RECT  0.125 -0.210 0.295 0.885 ;
        RECT  0.000 -0.210 0.125 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.980 2.310 8.400 2.730 ;
        RECT  7.720 2.035 7.980 2.730 ;
        RECT  7.245 2.310 7.720 2.730 ;
        RECT  6.985 2.015 7.245 2.730 ;
        RECT  5.415 2.310 6.985 2.730 ;
        RECT  5.155 2.260 5.415 2.730 ;
        RECT  3.405 2.310 5.155 2.730 ;
        RECT  3.145 2.220 3.405 2.730 ;
        RECT  2.820 2.310 3.145 2.730 ;
        RECT  2.560 2.220 2.820 2.730 ;
        RECT  1.560 2.310 2.560 2.730 ;
        RECT  1.440 1.995 1.560 2.730 ;
        RECT  0.295 2.310 1.440 2.730 ;
        RECT  0.125 1.930 0.295 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.400 2.520 ;
        LAYER M1 ;
        RECT  7.930 1.020 8.050 1.895 ;
        RECT  7.285 1.775 7.930 1.895 ;
        RECT  7.165 0.355 7.285 1.895 ;
        RECT  7.075 0.355 7.165 0.525 ;
        RECT  6.100 1.515 7.165 1.690 ;
        RECT  6.885 0.670 7.005 1.380 ;
        RECT  5.175 0.670 6.885 0.790 ;
        RECT  4.110 0.380 6.570 0.500 ;
        RECT  6.295 1.855 6.435 1.975 ;
        RECT  6.175 1.855 6.295 2.140 ;
        RECT  4.195 2.020 6.175 2.140 ;
        RECT  5.795 0.960 5.915 1.900 ;
        RECT  5.515 0.960 5.795 1.080 ;
        RECT  4.435 1.780 5.795 1.900 ;
        RECT  5.175 1.480 5.595 1.600 ;
        RECT  5.055 0.670 5.175 1.600 ;
        RECT  4.815 0.890 4.935 1.520 ;
        RECT  4.800 0.890 4.815 1.010 ;
        RECT  4.675 1.400 4.815 1.520 ;
        RECT  4.280 0.830 4.800 1.010 ;
        RECT  3.630 1.160 4.695 1.280 ;
        RECT  4.555 1.400 4.675 1.660 ;
        RECT  4.315 1.440 4.435 1.900 ;
        RECT  3.535 1.440 4.315 1.560 ;
        RECT  3.870 0.890 4.280 1.010 ;
        RECT  4.075 1.690 4.195 2.140 ;
        RECT  3.990 0.380 4.110 0.770 ;
        RECT  3.675 1.690 4.075 1.810 ;
        RECT  3.835 1.930 3.955 2.190 ;
        RECT  3.750 0.380 3.870 1.010 ;
        RECT  1.800 1.980 3.835 2.100 ;
        RECT  2.205 0.380 3.750 0.500 ;
        RECT  3.510 0.620 3.630 1.280 ;
        RECT  3.415 1.440 3.535 1.860 ;
        RECT  2.445 0.620 3.510 0.740 ;
        RECT  2.040 1.740 3.415 1.860 ;
        RECT  3.340 0.860 3.390 0.980 ;
        RECT  3.250 0.860 3.340 1.310 ;
        RECT  3.130 0.860 3.250 1.620 ;
        RECT  2.945 1.500 3.130 1.620 ;
        RECT  2.325 0.620 2.445 1.610 ;
        RECT  2.175 1.255 2.325 1.610 ;
        RECT  2.085 0.380 2.205 1.135 ;
        RECT  1.570 1.255 2.175 1.375 ;
        RECT  1.390 1.015 2.085 1.135 ;
        RECT  1.920 1.515 2.040 1.860 ;
        RECT  1.795 0.715 1.965 0.890 ;
        RECT  1.140 1.515 1.920 1.635 ;
        RECT  1.680 1.755 1.800 2.100 ;
        RECT  1.140 0.770 1.795 0.890 ;
        RECT  0.905 1.755 1.680 1.875 ;
        RECT  1.270 1.015 1.390 1.285 ;
        RECT  1.020 0.770 1.140 1.635 ;
        RECT  0.930 1.255 1.020 1.635 ;
        RECT  0.810 1.755 0.905 2.075 ;
        RECT  0.810 0.670 0.900 0.930 ;
        RECT  0.730 0.670 0.810 2.075 ;
        RECT  0.690 0.670 0.730 1.875 ;
    END
END DFFSRX2AD
MACRO DFFSRX4AD
    CLASS CORE ;
    FOREIGN DFFSRX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.120 1.925 8.445 2.185 ;
        END
        AntennaGateArea 0.15 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.880 3.010 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.030 0.415 9.170 1.655 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.930 1.005 10.010 1.515 ;
        RECT  9.770 0.415 9.930 1.985 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 1.185 0.535 1.615 ;
        END
        AntennaGateArea 0.065 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.565 0.990 2.730 1.540 ;
        END
        AntennaGateArea 0.119 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.275 -0.210 10.360 0.210 ;
        RECT  10.105 -0.210 10.275 0.810 ;
        RECT  9.555 -0.210 10.105 0.210 ;
        RECT  9.385 -0.210 9.555 0.810 ;
        RECT  8.835 -0.210 9.385 0.210 ;
        RECT  8.665 -0.210 8.835 0.415 ;
        RECT  7.900 -0.210 8.665 0.210 ;
        RECT  7.640 -0.210 7.900 0.590 ;
        RECT  2.885 -0.210 7.640 0.210 ;
        RECT  2.625 -0.210 2.885 0.260 ;
        RECT  1.585 -0.210 2.625 0.210 ;
        RECT  1.415 -0.210 1.585 0.650 ;
        RECT  0.295 -0.210 1.415 0.210 ;
        RECT  0.125 -0.210 0.295 0.850 ;
        RECT  0.000 -0.210 0.125 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.275 2.310 10.360 2.730 ;
        RECT  10.105 1.780 10.275 2.730 ;
        RECT  9.600 2.310 10.105 2.730 ;
        RECT  9.340 2.035 9.600 2.730 ;
        RECT  8.880 2.310 9.340 2.730 ;
        RECT  8.620 2.015 8.880 2.730 ;
        RECT  6.940 2.310 8.620 2.730 ;
        RECT  6.680 2.260 6.940 2.730 ;
        RECT  4.250 2.310 6.680 2.730 ;
        RECT  4.080 2.220 4.250 2.730 ;
        RECT  3.455 2.310 4.080 2.730 ;
        RECT  3.195 2.220 3.455 2.730 ;
        RECT  2.820 2.310 3.195 2.730 ;
        RECT  2.560 2.220 2.820 2.730 ;
        RECT  1.560 2.310 2.560 2.730 ;
        RECT  1.440 1.995 1.560 2.730 ;
        RECT  0.295 2.310 1.440 2.730 ;
        RECT  0.125 1.925 0.295 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.360 2.520 ;
        LAYER M1 ;
        RECT  9.530 1.020 9.650 1.895 ;
        RECT  8.910 1.775 9.530 1.895 ;
        RECT  8.790 0.720 8.910 1.895 ;
        RECT  8.310 0.720 8.790 0.840 ;
        RECT  7.665 1.540 8.790 1.725 ;
        RECT  8.460 1.045 8.630 1.215 ;
        RECT  7.100 1.070 8.460 1.190 ;
        RECT  8.160 0.370 8.300 0.490 ;
        RECT  8.040 0.370 8.160 0.830 ;
        RECT  7.495 0.710 8.040 0.830 ;
        RECT  7.830 1.890 8.000 2.010 ;
        RECT  7.710 1.890 7.830 2.140 ;
        RECT  5.480 2.020 7.710 2.140 ;
        RECT  7.375 0.530 7.495 0.830 ;
        RECT  7.360 1.510 7.480 1.860 ;
        RECT  7.325 0.530 7.375 0.765 ;
        RECT  6.830 1.740 7.360 1.860 ;
        RECT  7.220 0.530 7.325 0.650 ;
        RECT  7.100 1.500 7.240 1.620 ;
        RECT  7.100 0.380 7.220 0.650 ;
        RECT  4.670 0.380 7.100 0.500 ;
        RECT  6.980 0.770 7.100 1.620 ;
        RECT  6.910 0.770 6.980 0.890 ;
        RECT  6.650 0.620 6.910 0.890 ;
        RECT  6.710 1.010 6.830 1.860 ;
        RECT  6.550 1.010 6.710 1.130 ;
        RECT  5.105 1.740 6.710 1.860 ;
        RECT  6.430 0.770 6.650 0.890 ;
        RECT  6.310 0.620 6.430 1.620 ;
        RECT  5.550 0.620 6.310 0.740 ;
        RECT  5.940 1.500 6.310 1.620 ;
        RECT  5.820 0.860 6.190 0.980 ;
        RECT  5.700 0.860 5.820 1.620 ;
        RECT  5.030 0.860 5.700 0.980 ;
        RECT  5.560 1.500 5.700 1.620 ;
        RECT  5.460 1.100 5.580 1.360 ;
        RECT  5.220 1.980 5.480 2.140 ;
        RECT  3.755 1.160 5.460 1.280 ;
        RECT  4.730 2.020 5.220 2.140 ;
        RECT  4.985 1.440 5.105 1.860 ;
        RECT  4.770 0.810 5.030 0.980 ;
        RECT  3.495 1.440 4.985 1.560 ;
        RECT  4.240 0.860 4.770 0.980 ;
        RECT  4.610 1.690 4.730 2.140 ;
        RECT  4.550 0.380 4.670 0.740 ;
        RECT  3.655 1.690 4.610 1.810 ;
        RECT  4.410 0.620 4.550 0.740 ;
        RECT  4.370 1.930 4.490 2.190 ;
        RECT  1.800 1.980 4.370 2.100 ;
        RECT  4.120 0.380 4.240 0.980 ;
        RECT  2.205 0.380 4.120 0.500 ;
        RECT  3.635 0.620 3.755 1.280 ;
        RECT  2.445 0.620 3.635 0.740 ;
        RECT  3.375 1.440 3.495 1.860 ;
        RECT  3.340 0.860 3.390 0.980 ;
        RECT  2.050 1.740 3.375 1.860 ;
        RECT  3.250 0.860 3.340 1.310 ;
        RECT  3.130 0.860 3.250 1.620 ;
        RECT  2.945 1.500 3.130 1.620 ;
        RECT  2.325 0.620 2.445 1.610 ;
        RECT  2.175 1.255 2.325 1.610 ;
        RECT  2.085 0.380 2.205 1.135 ;
        RECT  1.570 1.255 2.175 1.375 ;
        RECT  1.390 1.015 2.085 1.135 ;
        RECT  1.930 1.515 2.050 1.860 ;
        RECT  1.795 0.715 1.965 0.890 ;
        RECT  1.140 1.515 1.930 1.635 ;
        RECT  1.680 1.755 1.800 2.100 ;
        RECT  1.140 0.770 1.795 0.890 ;
        RECT  0.905 1.755 1.680 1.875 ;
        RECT  1.270 1.015 1.390 1.285 ;
        RECT  1.020 0.770 1.140 1.635 ;
        RECT  0.930 1.255 1.020 1.635 ;
        RECT  0.810 1.755 0.905 2.075 ;
        RECT  0.810 0.670 0.900 0.930 ;
        RECT  0.730 0.670 0.810 2.075 ;
        RECT  0.690 0.670 0.730 1.875 ;
    END
END DFFSRX4AD
MACRO DFFSRXLAD
    CLASS CORE ;
    FOREIGN DFFSRXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.185 0.960 6.420 1.395 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.980 3.010 1.440 ;
        END
        AntennaGateArea 0.048 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.035 1.360 7.210 1.655 ;
        RECT  6.895 0.725 7.035 1.655 ;
        RECT  6.865 0.725 6.895 0.895 ;
        RECT  6.845 1.360 6.895 1.655 ;
        END
        AntennaDiffArea 0.143 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.610 0.690 7.770 1.700 ;
        END
        AntennaDiffArea 0.143 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.180 1.050 0.490 1.420 ;
        END
        AntennaGateArea 0.048 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.585 1.025 2.730 1.540 ;
        END
        AntennaGateArea 0.083 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.415 -0.210 7.840 0.210 ;
        RECT  7.245 -0.210 7.415 0.365 ;
        RECT  6.605 -0.210 7.245 0.210 ;
        RECT  6.435 -0.210 6.605 0.525 ;
        RECT  2.850 -0.210 6.435 0.210 ;
        RECT  2.590 -0.210 2.850 0.300 ;
        RECT  1.620 -0.210 2.590 0.210 ;
        RECT  1.450 -0.210 1.620 0.605 ;
        RECT  0.340 -0.210 1.450 0.210 ;
        RECT  0.170 -0.210 0.340 0.850 ;
        RECT  0.000 -0.210 0.170 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.420 2.310 7.840 2.730 ;
        RECT  7.160 2.015 7.420 2.730 ;
        RECT  6.945 2.310 7.160 2.730 ;
        RECT  6.685 2.015 6.945 2.730 ;
        RECT  5.020 2.310 6.685 2.730 ;
        RECT  4.760 2.210 5.020 2.730 ;
        RECT  3.480 2.310 4.760 2.730 ;
        RECT  3.220 2.040 3.480 2.730 ;
        RECT  2.820 2.310 3.220 2.730 ;
        RECT  2.560 2.075 2.820 2.730 ;
        RECT  1.560 2.310 2.560 2.730 ;
        RECT  1.440 1.995 1.560 2.730 ;
        RECT  0.340 2.310 1.440 2.730 ;
        RECT  0.170 1.685 0.340 2.730 ;
        RECT  0.000 2.310 0.170 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.840 2.520 ;
        LAYER M1 ;
        RECT  7.370 0.485 7.490 1.895 ;
        RECT  7.035 0.485 7.370 0.605 ;
        RECT  6.515 1.775 7.370 1.895 ;
        RECT  6.965 0.405 7.035 0.605 ;
        RECT  6.915 0.355 6.965 0.605 ;
        RECT  6.795 0.355 6.915 0.525 ;
        RECT  6.605 0.670 6.725 1.365 ;
        RECT  4.870 0.670 6.605 0.790 ;
        RECT  6.395 1.535 6.515 2.135 ;
        RECT  5.790 1.535 6.395 1.655 ;
        RECT  4.115 0.380 6.290 0.500 ;
        RECT  5.870 1.855 6.130 2.090 ;
        RECT  3.620 1.970 5.870 2.090 ;
        RECT  5.435 0.960 5.605 1.850 ;
        RECT  5.185 0.960 5.435 1.115 ;
        RECT  3.490 1.730 5.435 1.850 ;
        RECT  4.870 1.480 5.295 1.600 ;
        RECT  4.750 0.670 4.870 1.600 ;
        RECT  4.510 0.830 4.630 1.600 ;
        RECT  4.370 0.830 4.510 1.010 ;
        RECT  4.060 1.480 4.510 1.600 ;
        RECT  3.635 1.200 4.385 1.320 ;
        RECT  3.875 0.890 4.370 1.010 ;
        RECT  3.995 0.380 4.115 0.770 ;
        RECT  3.755 0.420 3.875 1.010 ;
        RECT  2.225 0.420 3.755 0.540 ;
        RECT  3.515 0.660 3.635 1.320 ;
        RECT  2.490 0.660 3.515 0.780 ;
        RECT  3.370 1.730 3.490 1.920 ;
        RECT  3.315 0.900 3.390 1.020 ;
        RECT  2.845 1.800 3.370 1.920 ;
        RECT  3.250 0.900 3.315 1.430 ;
        RECT  3.130 0.900 3.250 1.680 ;
        RECT  2.970 1.560 3.130 1.680 ;
        RECT  2.725 1.730 2.845 1.920 ;
        RECT  2.040 1.730 2.725 1.850 ;
        RECT  2.465 0.660 2.490 0.920 ;
        RECT  2.345 0.660 2.465 1.610 ;
        RECT  2.175 1.255 2.345 1.610 ;
        RECT  2.105 0.420 2.225 1.135 ;
        RECT  1.800 2.020 2.200 2.140 ;
        RECT  1.595 1.255 2.175 1.375 ;
        RECT  1.405 1.015 2.105 1.135 ;
        RECT  1.920 1.515 2.040 1.850 ;
        RECT  1.865 0.635 1.985 0.895 ;
        RECT  1.165 1.515 1.920 1.635 ;
        RECT  1.165 0.775 1.865 0.895 ;
        RECT  1.680 1.755 1.800 2.140 ;
        RECT  0.835 1.755 1.680 1.875 ;
        RECT  1.285 1.015 1.405 1.285 ;
        RECT  1.045 0.775 1.165 1.635 ;
        RECT  0.955 1.175 1.045 1.635 ;
        RECT  0.835 0.635 0.925 0.895 ;
        RECT  0.715 0.635 0.835 1.875 ;
    END
END DFFSRXLAD
MACRO DFFSX1AD
    CLASS CORE ;
    FOREIGN DFFSX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.510 1.100 4.690 1.620 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.270 0.690 5.370 0.950 ;
        RECT  5.270 1.330 5.370 1.590 ;
        RECT  5.110 0.690 5.270 1.590 ;
        END
        AntennaDiffArea 0.168 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.950 0.690 6.090 1.700 ;
        RECT  5.920 0.690 5.950 0.950 ;
        RECT  5.920 1.375 5.950 1.700 ;
        END
        AntennaDiffArea 0.203 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.510 1.440 ;
        RECT  0.260 1.180 0.350 1.440 ;
        END
        AntennaGateArea 0.077 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.525 0.910 2.775 1.090 ;
        RECT  2.405 0.910 2.525 1.275 ;
        END
        AntennaGateArea 0.089 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.865 -0.210 6.160 0.210 ;
        RECT  5.745 -0.210 5.865 0.430 ;
        RECT  4.840 -0.210 5.745 0.210 ;
        RECT  4.580 -0.210 4.840 0.300 ;
        RECT  2.605 -0.210 4.580 0.210 ;
        RECT  2.435 -0.210 2.605 0.370 ;
        RECT  1.335 -0.210 2.435 0.210 ;
        RECT  1.075 -0.210 1.335 0.300 ;
        RECT  0.295 -0.210 1.075 0.210 ;
        RECT  0.125 -0.210 0.295 0.385 ;
        RECT  0.000 -0.210 0.125 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.695 2.310 6.160 2.730 ;
        RECT  5.525 2.195 5.695 2.730 ;
        RECT  5.195 2.310 5.525 2.730 ;
        RECT  5.025 2.105 5.195 2.730 ;
        RECT  4.395 2.310 5.025 2.730 ;
        RECT  4.225 2.080 4.395 2.730 ;
        RECT  3.340 2.310 4.225 2.730 ;
        RECT  3.170 1.995 3.340 2.730 ;
        RECT  2.650 2.310 3.170 2.730 ;
        RECT  2.390 2.220 2.650 2.730 ;
        RECT  1.370 2.310 2.390 2.730 ;
        RECT  1.250 1.975 1.370 2.730 ;
        RECT  0.255 2.310 1.250 2.730 ;
        RECT  0.085 1.640 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.625 1.020 5.820 1.280 ;
        RECT  5.505 0.400 5.625 1.860 ;
        RECT  4.920 0.400 5.505 0.520 ;
        RECT  4.805 1.740 5.505 1.860 ;
        RECT  4.820 0.860 4.940 1.520 ;
        RECT  3.820 0.860 4.820 0.980 ;
        RECT  4.635 1.740 4.805 1.910 ;
        RECT  4.290 1.740 4.635 1.860 ;
        RECT  4.320 0.620 4.460 0.740 ;
        RECT  4.200 0.380 4.320 0.740 ;
        RECT  4.170 1.280 4.290 1.860 ;
        RECT  2.945 0.380 4.200 0.500 ;
        RECT  3.580 1.985 4.040 2.105 ;
        RECT  3.700 0.620 3.820 1.865 ;
        RECT  3.500 0.620 3.700 0.740 ;
        RECT  3.460 0.860 3.580 2.105 ;
        RECT  1.850 1.720 3.460 1.840 ;
        RECT  3.330 0.620 3.380 0.740 ;
        RECT  3.205 0.620 3.330 1.600 ;
        RECT  3.120 0.620 3.205 0.790 ;
        RECT  2.965 1.480 3.205 1.600 ;
        RECT  2.525 0.670 3.120 0.790 ;
        RECT  2.965 1.100 3.085 1.360 ;
        RECT  2.770 1.210 2.965 1.360 ;
        RECT  2.775 0.380 2.945 0.550 ;
        RECT  1.610 1.960 2.820 2.080 ;
        RECT  2.650 1.210 2.770 1.600 ;
        RECT  2.270 1.480 2.650 1.600 ;
        RECT  2.405 0.490 2.525 0.790 ;
        RECT  2.030 0.490 2.405 0.610 ;
        RECT  2.150 0.730 2.270 1.600 ;
        RECT  1.455 1.190 2.150 1.310 ;
        RECT  2.010 1.480 2.150 1.600 ;
        RECT  1.910 0.490 2.030 1.070 ;
        RECT  1.315 0.950 1.910 1.070 ;
        RECT  1.730 1.430 1.850 1.840 ;
        RECT  1.620 0.660 1.790 0.830 ;
        RECT  1.075 1.430 1.730 1.550 ;
        RECT  1.455 0.395 1.715 0.540 ;
        RECT  1.075 0.710 1.620 0.830 ;
        RECT  1.490 1.670 1.610 2.080 ;
        RECT  0.920 1.670 1.490 1.790 ;
        RECT  0.740 0.420 1.455 0.540 ;
        RECT  1.195 0.950 1.315 1.285 ;
        RECT  0.955 0.710 1.075 1.550 ;
        RECT  0.875 1.025 0.955 1.285 ;
        RECT  0.750 1.670 0.920 2.075 ;
        RECT  0.750 0.660 0.835 0.830 ;
        RECT  0.660 0.660 0.750 2.075 ;
        RECT  0.480 0.360 0.740 0.540 ;
        RECT  0.630 0.660 0.660 1.790 ;
    END
END DFFSX1AD
MACRO DFFSX2AD
    CLASS CORE ;
    FOREIGN DFFSX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.225 1.415 4.735 1.620 ;
        END
        AntennaGateArea 0.101 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.370 0.735 5.530 1.545 ;
        RECT  5.185 0.735 5.370 0.905 ;
        RECT  5.185 1.375 5.370 1.545 ;
        END
        AntennaDiffArea 0.287 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.950 0.380 6.090 1.895 ;
        RECT  5.920 0.380 5.950 0.900 ;
        RECT  5.920 1.375 5.950 1.895 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 1.130 0.310 1.390 ;
        RECT  0.070 0.865 0.240 1.390 ;
        END
        AntennaGateArea 0.077 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.910 2.775 1.090 ;
        RECT  2.330 0.910 2.450 1.275 ;
        END
        AntennaGateArea 0.096 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 -0.210 6.160 0.210 ;
        RECT  5.545 -0.210 5.715 0.535 ;
        RECT  4.620 -0.210 5.545 0.210 ;
        RECT  4.460 -0.210 4.620 0.735 ;
        RECT  2.620 -0.210 4.460 0.210 ;
        RECT  2.360 -0.210 2.620 0.260 ;
        RECT  1.275 -0.210 2.360 0.210 ;
        RECT  1.015 -0.210 1.275 0.240 ;
        RECT  0.255 -0.210 1.015 0.210 ;
        RECT  0.085 -0.210 0.255 0.360 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 2.310 6.160 2.730 ;
        RECT  5.545 1.980 5.715 2.730 ;
        RECT  5.085 2.310 5.545 2.730 ;
        RECT  4.915 2.225 5.085 2.730 ;
        RECT  4.345 2.310 4.915 2.730 ;
        RECT  4.175 2.080 4.345 2.730 ;
        RECT  3.270 2.310 4.175 2.730 ;
        RECT  3.100 2.020 3.270 2.730 ;
        RECT  2.610 2.310 3.100 2.730 ;
        RECT  2.350 2.220 2.610 2.730 ;
        RECT  1.330 2.310 2.350 2.730 ;
        RECT  1.210 2.010 1.330 2.730 ;
        RECT  0.255 2.310 1.210 2.730 ;
        RECT  0.085 1.615 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.800 1.000 5.830 1.260 ;
        RECT  5.680 1.000 5.800 1.860 ;
        RECT  5.060 1.740 5.680 1.860 ;
        RECT  4.940 0.350 5.060 1.860 ;
        RECT  4.765 1.740 4.940 1.860 ;
        RECT  4.765 1.000 4.820 1.260 ;
        RECT  4.645 0.860 4.765 1.260 ;
        RECT  4.595 1.740 4.765 1.910 ;
        RECT  3.760 0.860 4.645 0.980 ;
        RECT  4.040 1.740 4.595 1.860 ;
        RECT  4.160 0.620 4.310 0.740 ;
        RECT  4.040 1.175 4.190 1.295 ;
        RECT  4.040 0.380 4.160 0.740 ;
        RECT  2.960 0.380 4.040 0.500 ;
        RECT  3.920 1.175 4.040 1.860 ;
        RECT  3.510 1.985 4.010 2.105 ;
        RECT  3.640 0.620 3.760 1.735 ;
        RECT  3.440 0.620 3.640 0.740 ;
        RECT  3.390 0.860 3.510 2.105 ;
        RECT  1.810 1.710 3.390 1.830 ;
        RECT  3.260 0.620 3.320 0.740 ;
        RECT  3.140 0.620 3.260 1.590 ;
        RECT  3.060 0.620 3.140 0.790 ;
        RECT  2.935 1.470 3.140 1.590 ;
        RECT  2.515 0.670 3.060 0.790 ;
        RECT  2.900 1.090 3.020 1.350 ;
        RECT  2.700 0.380 2.960 0.540 ;
        RECT  2.710 1.230 2.900 1.350 ;
        RECT  1.570 1.960 2.790 2.080 ;
        RECT  2.590 1.230 2.710 1.590 ;
        RECT  2.210 1.470 2.590 1.590 ;
        RECT  2.395 0.380 2.515 0.790 ;
        RECT  1.970 0.380 2.395 0.500 ;
        RECT  2.090 0.620 2.210 1.590 ;
        RECT  1.970 1.235 2.090 1.590 ;
        RECT  1.850 0.380 1.970 1.115 ;
        RECT  1.500 1.235 1.970 1.355 ;
        RECT  1.345 0.995 1.850 1.115 ;
        RECT  1.690 1.480 1.810 1.830 ;
        RECT  1.560 0.620 1.730 0.790 ;
        RECT  1.050 1.480 1.690 1.600 ;
        RECT  1.515 0.350 1.655 0.470 ;
        RECT  1.450 1.720 1.570 2.080 ;
        RECT  1.050 0.670 1.560 0.790 ;
        RECT  1.395 0.350 1.515 0.500 ;
        RECT  0.865 1.720 1.450 1.840 ;
        RECT  0.735 0.380 1.395 0.500 ;
        RECT  1.225 0.995 1.345 1.335 ;
        RECT  1.175 1.165 1.225 1.335 ;
        RECT  0.930 0.670 1.050 1.600 ;
        RECT  0.815 1.025 0.930 1.285 ;
        RECT  0.695 1.720 0.865 1.915 ;
        RECT  0.690 0.620 0.810 0.790 ;
        RECT  0.475 0.350 0.735 0.500 ;
        RECT  0.690 1.720 0.695 1.840 ;
        RECT  0.570 0.620 0.690 1.840 ;
    END
END DFFSX2AD
MACRO DFFSX4AD
    CLASS CORE ;
    FOREIGN DFFSX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.045 1.470 5.575 1.610 ;
        RECT  4.875 1.440 5.045 1.610 ;
        END
        AntennaGateArea 0.146 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.945 0.380 6.115 1.620 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.995 6.930 1.515 ;
        RECT  6.690 0.380 6.850 1.985 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.130 0.490 1.655 ;
        RECT  0.215 1.130 0.350 1.390 ;
        END
        AntennaGateArea 0.084 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.500 0.900 2.775 1.095 ;
        RECT  2.380 0.900 2.500 1.160 ;
        END
        AntennaGateArea 0.113 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.195 -0.210 7.280 0.210 ;
        RECT  7.025 -0.210 7.195 0.830 ;
        RECT  6.475 -0.210 7.025 0.210 ;
        RECT  6.305 -0.210 6.475 0.830 ;
        RECT  5.755 -0.210 6.305 0.210 ;
        RECT  5.585 -0.210 5.755 0.415 ;
        RECT  5.165 -0.210 5.585 0.210 ;
        RECT  4.995 -0.210 5.165 0.415 ;
        RECT  2.770 -0.210 4.995 0.210 ;
        RECT  2.510 -0.210 2.770 0.260 ;
        RECT  1.425 -0.210 2.510 0.210 ;
        RECT  1.165 -0.210 1.425 0.415 ;
        RECT  0.260 -0.210 1.165 0.210 ;
        RECT  0.100 -0.210 0.260 0.915 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.195 2.310 7.280 2.730 ;
        RECT  7.025 1.645 7.195 2.730 ;
        RECT  6.475 2.310 7.025 2.730 ;
        RECT  6.305 2.030 6.475 2.730 ;
        RECT  5.755 2.310 6.305 2.730 ;
        RECT  5.585 2.030 5.755 2.730 ;
        RECT  4.935 2.310 5.585 2.730 ;
        RECT  4.765 2.065 4.935 2.730 ;
        RECT  3.695 2.310 4.765 2.730 ;
        RECT  3.525 2.065 3.695 2.730 ;
        RECT  3.290 2.310 3.525 2.730 ;
        RECT  3.120 2.065 3.290 2.730 ;
        RECT  2.660 2.310 3.120 2.730 ;
        RECT  2.400 1.965 2.660 2.730 ;
        RECT  1.350 2.310 2.400 2.730 ;
        RECT  1.190 2.025 1.350 2.730 ;
        RECT  0.265 2.310 1.190 2.730 ;
        RECT  0.095 1.790 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.280 2.520 ;
        LAYER M1 ;
        RECT  6.430 1.010 6.550 1.895 ;
        RECT  5.825 1.775 6.430 1.895 ;
        RECT  5.705 0.750 5.825 1.895 ;
        RECT  5.260 0.750 5.705 0.870 ;
        RECT  4.670 1.775 5.705 1.895 ;
        RECT  5.405 1.015 5.575 1.215 ;
        RECT  4.420 1.015 5.405 1.135 ;
        RECT  4.755 0.595 4.805 0.765 ;
        RECT  4.635 0.380 4.755 0.765 ;
        RECT  4.550 1.355 4.670 1.895 ;
        RECT  3.220 0.380 4.635 0.500 ;
        RECT  4.300 0.620 4.420 1.535 ;
        RECT  4.150 2.010 4.410 2.175 ;
        RECT  3.980 0.620 4.300 0.740 ;
        RECT  4.225 1.415 4.300 1.535 ;
        RECT  4.055 1.415 4.225 1.845 ;
        RECT  3.935 2.010 4.150 2.130 ;
        RECT  3.935 0.915 4.115 1.035 ;
        RECT  3.815 0.915 3.935 2.130 ;
        RECT  3.540 0.620 3.860 0.740 ;
        RECT  1.830 1.725 3.815 1.845 ;
        RECT  3.420 0.620 3.540 1.590 ;
        RECT  3.090 0.620 3.420 0.740 ;
        RECT  2.995 1.470 3.420 1.590 ;
        RECT  2.975 1.070 3.095 1.335 ;
        RECT  2.970 0.380 3.090 0.740 ;
        RECT  2.835 1.215 2.975 1.335 ;
        RECT  2.905 0.380 2.970 0.550 ;
        RECT  2.010 0.380 2.905 0.500 ;
        RECT  2.715 1.215 2.835 1.545 ;
        RECT  2.250 1.425 2.715 1.545 ;
        RECT  2.250 0.620 2.390 0.740 ;
        RECT  2.130 0.620 2.250 1.545 ;
        RECT  2.055 1.145 2.130 1.545 ;
        RECT  1.820 2.020 2.080 2.190 ;
        RECT  1.510 1.145 2.055 1.265 ;
        RECT  1.890 0.380 2.010 1.025 ;
        RECT  1.330 0.905 1.890 1.025 ;
        RECT  1.710 1.385 1.830 1.845 ;
        RECT  1.590 2.020 1.820 2.140 ;
        RECT  1.650 0.525 1.770 0.785 ;
        RECT  1.090 1.385 1.710 1.505 ;
        RECT  1.090 0.665 1.650 0.785 ;
        RECT  1.470 1.625 1.590 2.140 ;
        RECT  0.875 1.625 1.470 1.745 ;
        RECT  1.210 0.905 1.330 1.265 ;
        RECT  0.970 0.665 1.090 1.505 ;
        RECT  0.880 1.075 0.970 1.335 ;
        RECT  0.760 1.625 0.875 1.800 ;
        RECT  0.760 0.655 0.850 0.915 ;
        RECT  0.705 0.655 0.760 1.800 ;
        RECT  0.620 0.655 0.705 1.745 ;
    END
END DFFSX4AD
MACRO DFFSXLAD
    CLASS CORE ;
    FOREIGN DFFSXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.510 1.100 4.690 1.620 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.270 0.690 5.370 0.950 ;
        RECT  5.270 1.330 5.370 1.590 ;
        RECT  5.110 0.690 5.270 1.590 ;
        END
        AntennaDiffArea 0.124 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.950 0.690 6.090 1.700 ;
        RECT  5.920 0.690 5.950 0.950 ;
        RECT  5.920 1.375 5.950 1.700 ;
        END
        AntennaDiffArea 0.138 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.510 1.440 ;
        RECT  0.260 1.180 0.350 1.440 ;
        END
        AntennaGateArea 0.077 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.525 0.910 2.775 1.090 ;
        RECT  2.405 0.910 2.525 1.275 ;
        END
        AntennaGateArea 0.089 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.865 -0.210 6.160 0.210 ;
        RECT  5.745 -0.210 5.865 0.510 ;
        RECT  4.840 -0.210 5.745 0.210 ;
        RECT  4.580 -0.210 4.840 0.300 ;
        RECT  2.605 -0.210 4.580 0.210 ;
        RECT  2.435 -0.210 2.605 0.370 ;
        RECT  1.335 -0.210 2.435 0.210 ;
        RECT  1.075 -0.210 1.335 0.300 ;
        RECT  0.295 -0.210 1.075 0.210 ;
        RECT  0.125 -0.210 0.295 0.385 ;
        RECT  0.000 -0.210 0.125 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.695 2.310 6.160 2.730 ;
        RECT  5.525 2.005 5.695 2.730 ;
        RECT  5.195 2.310 5.525 2.730 ;
        RECT  5.025 1.980 5.195 2.730 ;
        RECT  4.395 2.310 5.025 2.730 ;
        RECT  4.225 2.080 4.395 2.730 ;
        RECT  3.340 2.310 4.225 2.730 ;
        RECT  3.170 1.995 3.340 2.730 ;
        RECT  2.650 2.310 3.170 2.730 ;
        RECT  2.390 2.220 2.650 2.730 ;
        RECT  1.370 2.310 2.390 2.730 ;
        RECT  1.250 1.975 1.370 2.730 ;
        RECT  0.255 2.310 1.250 2.730 ;
        RECT  0.085 1.640 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.625 1.020 5.820 1.280 ;
        RECT  5.505 0.400 5.625 1.860 ;
        RECT  4.920 0.400 5.505 0.520 ;
        RECT  4.805 1.740 5.505 1.860 ;
        RECT  4.820 0.860 4.940 1.520 ;
        RECT  3.820 0.860 4.820 0.980 ;
        RECT  4.635 1.740 4.805 1.910 ;
        RECT  4.290 1.740 4.635 1.860 ;
        RECT  4.320 0.620 4.460 0.740 ;
        RECT  4.200 0.380 4.320 0.740 ;
        RECT  4.170 1.280 4.290 1.860 ;
        RECT  2.945 0.380 4.200 0.500 ;
        RECT  3.580 1.985 4.040 2.105 ;
        RECT  3.700 0.620 3.820 1.865 ;
        RECT  3.500 0.620 3.700 0.740 ;
        RECT  3.460 0.860 3.580 2.105 ;
        RECT  1.850 1.720 3.460 1.840 ;
        RECT  3.330 0.620 3.380 0.740 ;
        RECT  3.205 0.620 3.330 1.600 ;
        RECT  3.120 0.620 3.205 0.790 ;
        RECT  2.965 1.480 3.205 1.600 ;
        RECT  2.525 0.670 3.120 0.790 ;
        RECT  2.965 1.100 3.085 1.360 ;
        RECT  2.770 1.210 2.965 1.360 ;
        RECT  2.775 0.380 2.945 0.550 ;
        RECT  1.610 1.960 2.820 2.080 ;
        RECT  2.650 1.210 2.770 1.600 ;
        RECT  2.270 1.480 2.650 1.600 ;
        RECT  2.405 0.490 2.525 0.790 ;
        RECT  2.030 0.490 2.405 0.610 ;
        RECT  2.150 0.730 2.270 1.600 ;
        RECT  1.455 1.190 2.150 1.310 ;
        RECT  2.010 1.480 2.150 1.600 ;
        RECT  1.910 0.490 2.030 1.070 ;
        RECT  1.315 0.950 1.910 1.070 ;
        RECT  1.730 1.430 1.850 1.840 ;
        RECT  1.620 0.660 1.790 0.830 ;
        RECT  1.075 1.430 1.730 1.550 ;
        RECT  1.455 0.395 1.715 0.540 ;
        RECT  1.075 0.710 1.620 0.830 ;
        RECT  1.490 1.670 1.610 2.080 ;
        RECT  0.920 1.670 1.490 1.790 ;
        RECT  0.740 0.420 1.455 0.540 ;
        RECT  1.195 0.950 1.315 1.285 ;
        RECT  0.955 0.710 1.075 1.550 ;
        RECT  0.875 1.025 0.955 1.285 ;
        RECT  0.750 1.670 0.920 2.075 ;
        RECT  0.750 0.660 0.835 0.830 ;
        RECT  0.660 0.660 0.750 2.075 ;
        RECT  0.480 0.360 0.740 0.540 ;
        RECT  0.630 0.660 0.660 1.790 ;
    END
END DFFSXLAD
MACRO DFFTRX1AD
    CLASS CORE ;
    FOREIGN DFFTRX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.585 1.095 0.950 ;
        END
        AntennaGateArea 0.043 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.330 1.140 5.530 1.380 ;
        RECT  5.170 0.660 5.330 1.590 ;
        END
        AntennaDiffArea 0.179 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.930 0.680 6.090 1.920 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 0.585 0.790 0.950 ;
        END
        AntennaGateArea 0.043 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.865 1.760 1.095 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 -0.210 6.160 0.210 ;
        RECT  5.545 -0.210 5.715 0.815 ;
        RECT  4.725 -0.210 5.545 0.210 ;
        RECT  4.465 -0.210 4.725 0.300 ;
        RECT  3.215 -0.210 4.465 0.210 ;
        RECT  2.955 -0.210 3.215 0.300 ;
        RECT  1.940 -0.210 2.955 0.210 ;
        RECT  1.680 -0.210 1.940 0.525 ;
        RECT  1.290 -0.210 1.680 0.210 ;
        RECT  1.030 -0.210 1.290 0.300 ;
        RECT  0.000 -0.210 1.030 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.740 2.310 6.160 2.730 ;
        RECT  5.480 2.220 5.740 2.730 ;
        RECT  4.810 2.310 5.480 2.730 ;
        RECT  4.550 2.240 4.810 2.730 ;
        RECT  3.230 2.310 4.550 2.730 ;
        RECT  3.205 1.830 3.230 2.730 ;
        RECT  3.085 1.780 3.205 2.730 ;
        RECT  3.060 1.830 3.085 2.730 ;
        RECT  1.940 2.310 3.060 2.730 ;
        RECT  1.680 2.220 1.940 2.730 ;
        RECT  1.040 2.310 1.680 2.730 ;
        RECT  0.780 2.215 1.040 2.730 ;
        RECT  0.000 2.310 0.780 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.690 1.010 5.810 1.895 ;
        RECT  5.040 1.765 5.690 1.895 ;
        RECT  4.920 0.540 5.040 2.100 ;
        RECT  4.860 0.540 4.920 0.800 ;
        RECT  4.860 1.715 4.920 2.100 ;
        RECT  4.430 1.980 4.860 2.100 ;
        RECT  4.680 1.025 4.800 1.545 ;
        RECT  4.555 0.850 4.680 1.850 ;
        RECT  4.105 0.850 4.555 0.970 ;
        RECT  3.735 1.730 4.555 1.850 ;
        RECT  4.260 1.980 4.430 2.185 ;
        RECT  3.955 1.175 4.215 1.575 ;
        RECT  3.905 0.540 4.105 0.970 ;
        RECT  3.785 1.175 3.955 1.300 ;
        RECT  3.665 0.420 3.785 1.300 ;
        RECT  2.710 0.420 3.665 0.540 ;
        RECT  3.545 1.450 3.615 1.970 ;
        RECT  3.425 0.660 3.545 1.970 ;
        RECT  3.390 0.660 3.425 0.920 ;
        RECT  3.035 0.800 3.390 0.920 ;
        RECT  3.185 1.040 3.305 1.605 ;
        RECT  2.660 1.485 3.185 1.605 ;
        RECT  2.915 0.800 3.035 1.365 ;
        RECT  2.775 1.245 2.915 1.365 ;
        RECT  2.280 0.380 2.710 0.540 ;
        RECT  2.630 0.740 2.660 0.860 ;
        RECT  2.630 1.485 2.660 2.095 ;
        RECT  2.510 0.740 2.630 2.095 ;
        RECT  2.400 0.740 2.510 0.860 ;
        RECT  2.430 1.780 2.510 2.095 ;
        RECT  0.255 1.975 2.430 2.095 ;
        RECT  2.250 0.380 2.280 1.600 ;
        RECT  2.160 0.380 2.250 1.740 ;
        RECT  2.075 0.380 2.160 0.525 ;
        RECT  2.130 1.480 2.160 1.740 ;
        RECT  0.495 1.480 2.130 1.600 ;
        RECT  1.920 0.645 2.040 1.360 ;
        RECT  1.350 1.240 1.920 1.360 ;
        RECT  1.350 0.575 1.505 0.745 ;
        RECT  0.400 1.735 1.380 1.855 ;
        RECT  1.230 0.575 1.350 1.360 ;
        RECT  0.470 1.125 1.230 1.245 ;
        RECT  0.325 1.390 0.495 1.600 ;
        RECT  0.350 0.985 0.470 1.245 ;
        RECT  0.205 0.425 0.315 0.595 ;
        RECT  0.205 1.720 0.255 2.095 ;
        RECT  0.085 0.425 0.205 2.095 ;
    END
END DFFTRX1AD
MACRO DFFTRX2AD
    CLASS CORE ;
    FOREIGN DFFTRX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.585 1.095 0.950 ;
        END
        AntennaGateArea 0.047 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.315 1.140 5.530 1.380 ;
        RECT  5.315 0.760 5.400 0.880 ;
        RECT  5.140 0.760 5.315 1.545 ;
        END
        AntennaDiffArea 0.322 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.680 6.090 2.020 ;
        RECT  5.930 0.365 6.050 2.020 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 0.585 0.790 0.950 ;
        END
        AntennaGateArea 0.058 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.865 1.755 1.095 ;
        END
        AntennaGateArea 0.08 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.760 -0.210 6.160 0.210 ;
        RECT  5.500 -0.210 5.760 0.390 ;
        RECT  4.745 -0.210 5.500 0.210 ;
        RECT  4.485 -0.210 4.745 0.300 ;
        RECT  3.215 -0.210 4.485 0.210 ;
        RECT  2.955 -0.210 3.215 0.260 ;
        RECT  1.940 -0.210 2.955 0.210 ;
        RECT  1.680 -0.210 1.940 0.525 ;
        RECT  1.290 -0.210 1.680 0.210 ;
        RECT  1.030 -0.210 1.290 0.355 ;
        RECT  0.000 -0.210 1.030 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.695 2.310 6.160 2.730 ;
        RECT  5.525 2.050 5.695 2.730 ;
        RECT  4.775 2.310 5.525 2.730 ;
        RECT  4.515 2.240 4.775 2.730 ;
        RECT  3.210 2.310 4.515 2.730 ;
        RECT  3.040 2.170 3.210 2.730 ;
        RECT  1.940 2.310 3.040 2.730 ;
        RECT  1.680 2.205 1.940 2.730 ;
        RECT  1.040 2.310 1.680 2.730 ;
        RECT  0.780 2.205 1.040 2.730 ;
        RECT  0.000 2.310 0.780 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.690 0.520 5.810 1.930 ;
        RECT  4.980 0.520 5.690 0.640 ;
        RECT  5.035 1.810 5.690 1.930 ;
        RECT  4.865 1.775 5.035 1.950 ;
        RECT  4.860 0.520 4.980 0.800 ;
        RECT  4.445 1.830 4.865 1.950 ;
        RECT  4.710 0.940 4.830 1.460 ;
        RECT  4.505 1.085 4.710 1.205 ;
        RECT  4.385 0.845 4.505 1.710 ;
        RECT  4.325 1.830 4.445 2.090 ;
        RECT  4.045 0.845 4.385 0.965 ;
        RECT  3.735 1.590 4.385 1.710 ;
        RECT  3.955 1.175 4.215 1.430 ;
        RECT  3.785 2.070 4.185 2.190 ;
        RECT  3.925 0.540 4.045 0.965 ;
        RECT  3.785 1.175 3.955 1.300 ;
        RECT  3.665 0.380 3.785 1.300 ;
        RECT  3.665 1.930 3.785 2.190 ;
        RECT  2.710 0.380 3.665 0.500 ;
        RECT  2.755 1.930 3.665 2.050 ;
        RECT  3.545 1.450 3.615 1.710 ;
        RECT  3.425 0.620 3.545 1.710 ;
        RECT  3.380 0.620 3.425 0.910 ;
        RECT  3.035 0.790 3.380 0.910 ;
        RECT  3.185 1.030 3.305 1.810 ;
        RECT  2.515 1.690 3.185 1.810 ;
        RECT  2.915 0.790 3.035 1.290 ;
        RECT  2.775 1.170 2.915 1.290 ;
        RECT  2.635 1.930 2.755 2.190 ;
        RECT  2.275 0.380 2.710 0.530 ;
        RECT  2.515 0.690 2.660 0.810 ;
        RECT  2.395 0.690 2.515 2.085 ;
        RECT  0.255 1.965 2.395 2.085 ;
        RECT  2.155 0.380 2.275 1.635 ;
        RECT  2.075 0.380 2.155 0.530 ;
        RECT  2.105 1.465 2.155 1.635 ;
        RECT  0.495 1.465 2.105 1.585 ;
        RECT  1.915 0.775 2.035 1.345 ;
        RECT  1.350 1.225 1.915 1.345 ;
        RECT  1.350 0.560 1.505 0.730 ;
        RECT  0.400 1.725 1.380 1.845 ;
        RECT  1.230 0.560 1.350 1.345 ;
        RECT  0.470 1.125 1.230 1.245 ;
        RECT  0.325 1.390 0.495 1.585 ;
        RECT  0.350 0.985 0.470 1.245 ;
        RECT  0.205 0.425 0.315 0.595 ;
        RECT  0.205 1.720 0.255 2.085 ;
        RECT  0.085 0.425 0.205 2.085 ;
    END
END DFFTRX2AD
MACRO DFFTRX4AD
    CLASS CORE ;
    FOREIGN DFFTRX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.585 1.095 0.950 ;
        RECT  0.930 0.585 1.050 1.090 ;
        RECT  0.910 0.585 0.930 0.950 ;
        END
        AntennaGateArea 0.08 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.785 0.405 6.955 1.555 ;
        RECT  6.715 1.005 6.785 1.555 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.695 1.005 7.770 1.515 ;
        RECT  7.505 0.405 7.695 1.945 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.585 0.790 0.950 ;
        RECT  0.630 0.585 0.750 1.090 ;
        RECT  0.600 0.585 0.630 0.950 ;
        END
        AntennaGateArea 0.109 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.865 1.755 1.095 ;
        END
        AntennaGateArea 0.119 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.010 -0.210 8.120 0.210 ;
        RECT  7.890 -0.210 8.010 0.815 ;
        RECT  7.315 -0.210 7.890 0.210 ;
        RECT  7.145 -0.210 7.315 0.770 ;
        RECT  6.570 -0.210 7.145 0.210 ;
        RECT  6.450 -0.210 6.570 0.810 ;
        RECT  5.910 -0.210 6.450 0.210 ;
        RECT  5.650 -0.210 5.910 0.855 ;
        RECT  4.055 -0.210 5.650 0.210 ;
        RECT  3.795 -0.210 4.055 0.260 ;
        RECT  3.295 -0.210 3.795 0.210 ;
        RECT  3.035 -0.210 3.295 0.260 ;
        RECT  1.940 -0.210 3.035 0.210 ;
        RECT  1.680 -0.210 1.940 0.525 ;
        RECT  1.290 -0.210 1.680 0.210 ;
        RECT  1.030 -0.210 1.290 0.330 ;
        RECT  0.000 -0.210 1.030 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.010 2.310 8.120 2.730 ;
        RECT  7.890 1.665 8.010 2.730 ;
        RECT  7.315 2.310 7.890 2.730 ;
        RECT  7.145 1.975 7.315 2.730 ;
        RECT  6.570 2.310 7.145 2.730 ;
        RECT  6.450 1.960 6.570 2.730 ;
        RECT  5.870 2.310 6.450 2.730 ;
        RECT  5.700 2.160 5.870 2.730 ;
        RECT  3.925 2.310 5.700 2.730 ;
        RECT  3.805 2.170 3.925 2.730 ;
        RECT  3.160 2.310 3.805 2.730 ;
        RECT  2.990 2.170 3.160 2.730 ;
        RECT  2.030 2.310 2.990 2.730 ;
        RECT  1.770 2.190 2.030 2.730 ;
        RECT  1.070 2.310 1.770 2.730 ;
        RECT  0.810 2.260 1.070 2.730 ;
        RECT  0.000 2.310 0.810 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.120 2.520 ;
        LAYER M1 ;
        RECT  7.335 1.010 7.385 1.270 ;
        RECT  7.215 1.010 7.335 1.810 ;
        RECT  6.330 1.680 7.215 1.810 ;
        RECT  6.250 0.620 6.330 2.040 ;
        RECT  6.205 0.620 6.250 2.070 ;
        RECT  6.100 0.620 6.205 0.880 ;
        RECT  6.080 1.640 6.205 2.070 ;
        RECT  5.450 1.920 6.080 2.040 ;
        RECT  5.680 1.000 6.015 1.520 ;
        RECT  5.560 0.975 5.680 1.760 ;
        RECT  5.160 0.975 5.560 1.095 ;
        RECT  5.090 1.640 5.560 1.760 ;
        RECT  5.260 1.340 5.400 1.460 ;
        RECT  5.140 1.215 5.260 1.460 ;
        RECT  5.040 0.650 5.160 1.095 ;
        RECT  4.880 1.215 5.140 1.335 ;
        RECT  4.970 1.640 5.090 1.900 ;
        RECT  4.445 1.780 4.970 1.900 ;
        RECT  4.760 0.380 4.880 1.335 ;
        RECT  4.590 1.455 4.850 1.640 ;
        RECT  2.710 0.380 4.760 0.500 ;
        RECT  4.280 1.215 4.760 1.335 ;
        RECT  3.605 0.690 4.610 0.810 ;
        RECT  3.605 1.455 4.590 1.575 ;
        RECT  4.325 1.695 4.445 1.900 ;
        RECT  4.275 1.695 4.325 1.865 ;
        RECT  4.160 0.940 4.280 1.335 ;
        RECT  4.045 1.930 4.165 2.190 ;
        RECT  2.755 1.930 4.045 2.050 ;
        RECT  3.545 0.690 3.605 1.575 ;
        RECT  3.485 0.690 3.545 1.715 ;
        RECT  3.000 0.690 3.485 0.810 ;
        RECT  3.425 1.455 3.485 1.715 ;
        RECT  3.185 1.030 3.305 1.810 ;
        RECT  2.515 1.690 3.185 1.810 ;
        RECT  3.000 1.170 3.035 1.290 ;
        RECT  2.880 0.690 3.000 1.290 ;
        RECT  2.775 1.170 2.880 1.290 ;
        RECT  2.635 1.930 2.755 2.190 ;
        RECT  2.275 0.380 2.710 0.530 ;
        RECT  2.515 0.690 2.660 0.810 ;
        RECT  2.395 0.690 2.515 2.010 ;
        RECT  1.620 1.890 2.395 2.010 ;
        RECT  2.155 0.380 2.275 1.740 ;
        RECT  2.075 0.380 2.155 0.530 ;
        RECT  2.105 1.540 2.155 1.740 ;
        RECT  1.250 1.540 2.105 1.660 ;
        RECT  1.915 0.985 2.035 1.420 ;
        RECT  1.490 1.300 1.915 1.420 ;
        RECT  1.500 1.890 1.620 2.140 ;
        RECT  1.350 0.575 1.505 0.745 ;
        RECT  0.285 2.020 1.500 2.140 ;
        RECT  1.370 1.220 1.490 1.420 ;
        RECT  0.645 1.780 1.380 1.900 ;
        RECT  1.350 1.220 1.370 1.340 ;
        RECT  1.230 0.575 1.350 1.340 ;
        RECT  1.130 1.460 1.250 1.660 ;
        RECT  0.430 1.220 1.230 1.340 ;
        RECT  0.310 1.460 1.130 1.580 ;
        RECT  0.475 1.730 0.645 1.900 ;
        RECT  0.310 1.080 0.430 1.340 ;
        RECT  0.190 0.330 0.360 0.710 ;
        RECT  0.190 1.710 0.285 2.140 ;
        RECT  0.115 0.330 0.190 2.140 ;
        RECT  0.100 0.330 0.115 1.855 ;
        RECT  0.070 0.565 0.100 1.855 ;
    END
END DFFTRX4AD
MACRO DFFTRXLAD
    CLASS CORE ;
    FOREIGN DFFTRXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.585 1.095 0.950 ;
        END
        AntennaGateArea 0.043 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.125 1.140 5.250 1.380 ;
        RECT  4.955 0.735 5.125 1.545 ;
        END
        AntennaDiffArea 0.143 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.670 0.680 5.810 1.655 ;
        RECT  5.650 0.680 5.670 0.940 ;
        RECT  5.650 1.395 5.670 1.655 ;
        END
        AntennaDiffArea 0.143 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 0.585 0.790 0.950 ;
        END
        AntennaGateArea 0.043 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.865 1.760 1.095 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.550 -0.210 5.880 0.210 ;
        RECT  5.290 -0.210 5.550 0.375 ;
        RECT  4.670 -0.210 5.290 0.210 ;
        RECT  4.410 -0.210 4.670 0.295 ;
        RECT  3.215 -0.210 4.410 0.210 ;
        RECT  2.955 -0.210 3.215 0.300 ;
        RECT  1.940 -0.210 2.955 0.210 ;
        RECT  1.680 -0.210 1.940 0.525 ;
        RECT  1.290 -0.210 1.680 0.210 ;
        RECT  1.030 -0.210 1.290 0.300 ;
        RECT  0.000 -0.210 1.030 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.460 2.310 5.880 2.730 ;
        RECT  5.200 2.030 5.460 2.730 ;
        RECT  4.700 2.310 5.200 2.730 ;
        RECT  4.440 1.905 4.700 2.730 ;
        RECT  3.230 2.310 4.440 2.730 ;
        RECT  3.205 1.830 3.230 2.730 ;
        RECT  3.085 1.780 3.205 2.730 ;
        RECT  3.060 1.830 3.085 2.730 ;
        RECT  1.940 2.310 3.060 2.730 ;
        RECT  1.680 2.220 1.940 2.730 ;
        RECT  1.040 2.310 1.680 2.730 ;
        RECT  0.780 2.215 1.040 2.730 ;
        RECT  0.000 2.310 0.780 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.880 2.520 ;
        LAYER M1 ;
        RECT  5.530 1.010 5.550 1.270 ;
        RECT  5.410 0.495 5.530 1.785 ;
        RECT  5.005 0.495 5.410 0.615 ;
        RECT  5.010 1.665 5.410 1.785 ;
        RECT  4.890 1.665 5.010 2.130 ;
        RECT  4.835 0.375 5.005 0.615 ;
        RECT  4.495 1.665 4.890 1.785 ;
        RECT  4.710 0.885 4.830 1.405 ;
        RECT  4.255 1.085 4.710 1.205 ;
        RECT  4.375 1.350 4.495 1.785 ;
        RECT  4.135 0.850 4.255 1.850 ;
        RECT  4.025 0.850 4.135 0.970 ;
        RECT  3.735 1.730 4.135 1.850 ;
        RECT  3.905 0.540 4.025 0.970 ;
        RECT  3.895 1.225 4.015 1.610 ;
        RECT  3.785 1.225 3.895 1.345 ;
        RECT  3.665 0.330 3.785 1.345 ;
        RECT  3.525 0.330 3.665 0.540 ;
        RECT  3.545 1.735 3.590 1.905 ;
        RECT  3.425 0.660 3.545 1.905 ;
        RECT  2.710 0.420 3.525 0.540 ;
        RECT  3.390 0.660 3.425 0.920 ;
        RECT  3.420 1.735 3.425 1.905 ;
        RECT  3.035 0.800 3.390 0.920 ;
        RECT  3.185 1.040 3.305 1.605 ;
        RECT  2.660 1.485 3.185 1.605 ;
        RECT  2.915 0.800 3.035 1.365 ;
        RECT  2.775 1.245 2.915 1.365 ;
        RECT  2.280 0.380 2.710 0.540 ;
        RECT  2.630 0.740 2.660 0.860 ;
        RECT  2.630 1.485 2.660 2.095 ;
        RECT  2.510 0.740 2.630 2.095 ;
        RECT  2.400 0.740 2.510 0.860 ;
        RECT  2.430 1.780 2.510 2.095 ;
        RECT  0.255 1.975 2.430 2.095 ;
        RECT  2.250 0.380 2.280 1.600 ;
        RECT  2.160 0.380 2.250 1.740 ;
        RECT  2.075 0.380 2.160 0.525 ;
        RECT  2.130 1.480 2.160 1.740 ;
        RECT  0.495 1.480 2.130 1.600 ;
        RECT  1.920 0.645 2.040 1.360 ;
        RECT  1.350 1.240 1.920 1.360 ;
        RECT  1.350 0.575 1.505 0.745 ;
        RECT  0.400 1.735 1.380 1.855 ;
        RECT  1.230 0.575 1.350 1.360 ;
        RECT  0.470 1.125 1.230 1.245 ;
        RECT  0.325 1.390 0.495 1.600 ;
        RECT  0.350 0.985 0.470 1.245 ;
        RECT  0.205 0.425 0.315 0.595 ;
        RECT  0.205 1.720 0.255 2.095 ;
        RECT  0.085 0.425 0.205 2.095 ;
    END
END DFFTRXLAD
MACRO DFFX1AD
    CLASS CORE ;
    FOREIGN DFFX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.950 0.700 6.090 1.770 ;
        RECT  5.905 0.700 5.950 0.870 ;
        RECT  5.930 1.470 5.950 1.770 ;
        END
        AntennaDiffArea 0.207 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 0.755 5.530 1.480 ;
        RECT  5.365 0.755 5.390 0.895 ;
        RECT  5.280 1.340 5.390 1.480 ;
        RECT  5.195 0.725 5.365 0.895 ;
        RECT  5.160 1.340 5.280 1.600 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.740 0.235 1.380 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.705 1.190 1.935 1.610 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.790 -0.210 6.160 0.210 ;
        RECT  5.530 -0.210 5.790 0.380 ;
        RECT  4.635 -0.210 5.530 0.210 ;
        RECT  4.465 -0.210 4.635 0.325 ;
        RECT  3.480 -0.210 4.465 0.210 ;
        RECT  3.220 -0.210 3.480 0.300 ;
        RECT  2.520 -0.210 3.220 0.210 ;
        RECT  2.260 -0.210 2.520 0.300 ;
        RECT  1.790 -0.210 2.260 0.210 ;
        RECT  1.530 -0.210 1.790 0.300 ;
        RECT  0.265 -0.210 1.530 0.210 ;
        RECT  0.095 -0.210 0.265 0.535 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.730 2.310 6.160 2.730 ;
        RECT  5.470 2.020 5.730 2.730 ;
        RECT  4.670 2.310 5.470 2.730 ;
        RECT  4.410 2.060 4.670 2.730 ;
        RECT  3.280 2.310 4.410 2.730 ;
        RECT  3.020 2.220 3.280 2.730 ;
        RECT  2.230 2.310 3.020 2.730 ;
        RECT  1.970 2.220 2.230 2.730 ;
        RECT  1.500 2.310 1.970 2.730 ;
        RECT  1.240 2.220 1.500 2.730 ;
        RECT  0.240 2.310 1.240 2.730 ;
        RECT  0.120 1.550 0.240 2.730 ;
        RECT  0.000 2.310 0.120 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.810 1.010 5.830 1.270 ;
        RECT  5.690 1.010 5.810 1.840 ;
        RECT  5.040 1.720 5.690 1.840 ;
        RECT  4.940 0.595 5.040 1.840 ;
        RECT  4.920 0.595 4.940 1.940 ;
        RECT  4.845 0.595 4.920 0.765 ;
        RECT  4.820 1.505 4.920 1.940 ;
        RECT  4.140 1.820 4.820 1.940 ;
        RECT  4.530 1.000 4.790 1.260 ;
        RECT  4.410 0.690 4.530 1.670 ;
        RECT  4.040 0.690 4.410 0.810 ;
        RECT  3.850 1.550 4.410 1.670 ;
        RECT  4.130 0.940 4.260 1.060 ;
        RECT  4.000 0.940 4.130 1.430 ;
        RECT  3.920 0.550 4.040 0.810 ;
        RECT  3.510 1.310 4.000 1.430 ;
        RECT  3.775 0.930 3.880 1.190 ;
        RECT  3.730 1.550 3.850 1.820 ;
        RECT  3.510 1.980 3.800 2.100 ;
        RECT  3.655 0.420 3.775 1.190 ;
        RECT  3.090 0.420 3.655 0.540 ;
        RECT  3.390 0.800 3.510 2.100 ;
        RECT  3.240 0.800 3.390 0.920 ;
        RECT  0.590 1.980 3.390 2.100 ;
        RECT  3.150 1.100 3.270 1.860 ;
        RECT  3.120 0.660 3.240 0.920 ;
        RECT  2.490 1.740 3.150 1.860 ;
        RECT  3.000 0.380 3.090 0.540 ;
        RECT  2.880 0.380 3.000 1.620 ;
        RECT  2.830 0.380 2.880 0.540 ;
        RECT  2.630 1.500 2.880 1.620 ;
        RECT  2.430 0.420 2.830 0.540 ;
        RECT  2.640 0.660 2.760 1.325 ;
        RECT  2.490 1.205 2.640 1.325 ;
        RECT  2.370 1.205 2.490 1.860 ;
        RECT  2.310 0.420 2.430 0.830 ;
        RECT  1.420 1.740 2.370 1.860 ;
        RECT  1.230 0.710 2.310 0.830 ;
        RECT  2.110 0.950 2.230 1.230 ;
        RECT  1.955 0.365 2.125 0.540 ;
        RECT  1.475 0.950 2.110 1.070 ;
        RECT  0.710 0.420 1.955 0.540 ;
        RECT  1.355 0.950 1.475 1.160 ;
        RECT  1.290 1.290 1.420 1.860 ;
        RECT  0.970 1.040 1.355 1.160 ;
        RECT  1.160 1.290 1.290 1.410 ;
        RECT  1.110 0.660 1.230 0.920 ;
        RECT  0.860 0.660 0.970 1.160 ;
        RECT  0.850 0.660 0.860 1.770 ;
        RECT  0.740 1.040 0.850 1.770 ;
        RECT  0.590 0.420 0.710 0.900 ;
        RECT  0.470 0.680 0.590 2.100 ;
    END
END DFFX1AD
MACRO DFFX2AD
    CLASS CORE ;
    FOREIGN DFFX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 0.865 6.090 1.375 ;
        RECT  5.930 0.420 6.050 2.010 ;
        END
        AntennaDiffArea 0.373 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 0.760 5.530 1.515 ;
        RECT  5.140 0.760 5.390 0.900 ;
        RECT  5.355 1.375 5.390 1.515 ;
        RECT  5.185 1.375 5.355 1.545 ;
        END
        AntennaDiffArea 0.353 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.760 0.235 1.375 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.705 1.190 1.935 1.610 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.760 -0.210 6.160 0.210 ;
        RECT  5.500 -0.210 5.760 0.390 ;
        RECT  4.600 -0.210 5.500 0.210 ;
        RECT  4.480 -0.210 4.600 0.370 ;
        RECT  3.410 -0.210 4.480 0.210 ;
        RECT  3.150 -0.210 3.410 0.300 ;
        RECT  2.460 -0.210 3.150 0.210 ;
        RECT  2.200 -0.210 2.460 0.300 ;
        RECT  1.740 -0.210 2.200 0.210 ;
        RECT  1.480 -0.210 1.740 0.300 ;
        RECT  0.230 -0.210 1.480 0.210 ;
        RECT  0.110 -0.210 0.230 0.580 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.760 2.310 6.160 2.730 ;
        RECT  5.500 2.010 5.760 2.730 ;
        RECT  4.635 2.310 5.500 2.730 ;
        RECT  4.375 2.060 4.635 2.730 ;
        RECT  3.210 2.310 4.375 2.730 ;
        RECT  2.950 2.220 3.210 2.730 ;
        RECT  2.190 2.310 2.950 2.730 ;
        RECT  1.930 2.220 2.190 2.730 ;
        RECT  1.460 2.310 1.930 2.730 ;
        RECT  1.200 2.220 1.460 2.730 ;
        RECT  0.230 2.310 1.200 2.730 ;
        RECT  0.110 1.550 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.690 0.520 5.810 1.830 ;
        RECT  5.055 0.520 5.690 0.640 ;
        RECT  4.970 1.710 5.690 1.830 ;
        RECT  4.530 1.045 5.135 1.215 ;
        RECT  4.885 0.385 5.055 0.640 ;
        RECT  4.850 1.445 4.970 1.940 ;
        RECT  4.080 1.820 4.850 1.940 ;
        RECT  4.410 0.690 4.530 1.670 ;
        RECT  3.970 0.690 4.410 0.810 ;
        RECT  3.780 1.550 4.410 1.670 ;
        RECT  4.050 0.940 4.190 1.060 ;
        RECT  3.930 0.940 4.050 1.430 ;
        RECT  3.945 2.070 4.040 2.190 ;
        RECT  3.850 0.550 3.970 0.810 ;
        RECT  3.780 1.980 3.945 2.190 ;
        RECT  3.440 1.310 3.930 1.430 ;
        RECT  3.680 0.930 3.810 1.190 ;
        RECT  3.660 1.550 3.780 1.830 ;
        RECT  3.440 1.980 3.780 2.100 ;
        RECT  3.560 0.420 3.680 1.190 ;
        RECT  3.020 0.420 3.560 0.540 ;
        RECT  3.320 0.800 3.440 2.100 ;
        RECT  3.170 0.800 3.320 0.920 ;
        RECT  0.590 1.980 3.320 2.100 ;
        RECT  3.080 1.100 3.200 1.860 ;
        RECT  3.050 0.660 3.170 0.920 ;
        RECT  2.430 1.740 3.080 1.860 ;
        RECT  2.930 0.380 3.020 0.540 ;
        RECT  2.810 0.380 2.930 1.620 ;
        RECT  2.760 0.380 2.810 0.540 ;
        RECT  2.560 1.500 2.810 1.620 ;
        RECT  2.410 0.420 2.760 0.540 ;
        RECT  2.570 0.660 2.690 1.325 ;
        RECT  2.430 1.205 2.570 1.325 ;
        RECT  2.310 1.205 2.430 1.860 ;
        RECT  2.290 0.420 2.410 0.830 ;
        RECT  1.535 1.740 2.310 1.860 ;
        RECT  1.200 0.710 2.290 0.830 ;
        RECT  2.070 0.950 2.190 1.230 ;
        RECT  1.905 0.365 2.075 0.540 ;
        RECT  1.440 0.950 2.070 1.070 ;
        RECT  0.680 0.420 1.905 0.540 ;
        RECT  1.415 1.290 1.535 1.860 ;
        RECT  1.320 0.950 1.440 1.160 ;
        RECT  1.140 1.290 1.415 1.410 ;
        RECT  0.940 1.040 1.320 1.160 ;
        RECT  1.080 0.660 1.200 0.920 ;
        RECT  0.840 0.660 0.940 1.160 ;
        RECT  0.820 0.660 0.840 1.805 ;
        RECT  0.720 1.040 0.820 1.805 ;
        RECT  0.590 0.420 0.680 0.900 ;
        RECT  0.560 0.420 0.590 2.100 ;
        RECT  0.470 0.680 0.560 2.100 ;
    END
END DFFX2AD
MACRO DFFX4AD
    CLASS CORE ;
    FOREIGN DFFX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.430 1.005 7.490 1.515 ;
        RECT  7.410 0.430 7.430 1.515 ;
        RECT  7.250 0.430 7.410 2.120 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.510 0.430 6.650 1.590 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.765 0.235 1.375 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.935 1.190 1.990 1.310 ;
        RECT  1.705 1.190 1.935 1.610 ;
        END
        AntennaGateArea 0.095 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.755 -0.210 7.840 0.210 ;
        RECT  7.585 -0.210 7.755 0.830 ;
        RECT  7.035 -0.210 7.585 0.210 ;
        RECT  6.865 -0.210 7.035 0.785 ;
        RECT  6.315 -0.210 6.865 0.210 ;
        RECT  6.145 -0.210 6.315 0.530 ;
        RECT  5.730 -0.210 6.145 0.210 ;
        RECT  5.470 -0.210 5.730 0.300 ;
        RECT  4.840 -0.210 5.470 0.210 ;
        RECT  4.580 -0.210 4.840 0.300 ;
        RECT  3.580 -0.210 4.580 0.210 ;
        RECT  3.320 -0.210 3.580 0.300 ;
        RECT  2.520 -0.210 3.320 0.210 ;
        RECT  2.260 -0.210 2.520 0.300 ;
        RECT  1.800 -0.210 2.260 0.210 ;
        RECT  1.540 -0.210 1.800 0.300 ;
        RECT  0.265 -0.210 1.540 0.210 ;
        RECT  0.095 -0.210 0.265 0.525 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.730 2.310 7.840 2.730 ;
        RECT  7.610 1.550 7.730 2.730 ;
        RECT  7.080 2.310 7.610 2.730 ;
        RECT  6.820 2.005 7.080 2.730 ;
        RECT  6.360 2.310 6.820 2.730 ;
        RECT  6.100 2.010 6.360 2.730 ;
        RECT  5.630 2.310 6.100 2.730 ;
        RECT  5.370 2.030 5.630 2.730 ;
        RECT  4.540 2.310 5.370 2.730 ;
        RECT  4.280 1.785 4.540 2.730 ;
        RECT  3.290 2.310 4.280 2.730 ;
        RECT  3.030 2.220 3.290 2.730 ;
        RECT  2.220 2.310 3.030 2.730 ;
        RECT  1.960 2.220 2.220 2.730 ;
        RECT  1.500 2.310 1.960 2.730 ;
        RECT  1.240 2.220 1.500 2.730 ;
        RECT  0.265 2.310 1.240 2.730 ;
        RECT  0.095 1.585 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.840 2.520 ;
        LAYER M1 ;
        RECT  7.010 1.020 7.130 1.875 ;
        RECT  6.390 1.755 7.010 1.875 ;
        RECT  6.270 0.680 6.390 1.875 ;
        RECT  5.760 0.680 6.270 0.800 ;
        RECT  5.975 1.755 6.270 1.875 ;
        RECT  5.580 1.000 6.090 1.260 ;
        RECT  5.805 1.440 5.975 1.875 ;
        RECT  5.340 1.755 5.805 1.875 ;
        RECT  5.460 0.520 5.580 1.585 ;
        RECT  4.140 0.520 5.460 0.640 ;
        RECT  3.930 1.465 5.460 1.585 ;
        RECT  5.080 1.755 5.340 1.905 ;
        RECT  5.070 0.760 5.190 1.345 ;
        RECT  3.550 1.225 5.070 1.345 ;
        RECT  4.770 0.845 4.890 1.105 ;
        RECT  3.900 0.845 4.770 0.990 ;
        RECT  4.020 0.370 4.140 0.640 ;
        RECT  3.550 1.980 4.060 2.190 ;
        RECT  3.670 1.465 3.930 1.735 ;
        RECT  3.780 0.420 3.900 0.990 ;
        RECT  3.050 0.420 3.780 0.540 ;
        RECT  3.540 0.800 3.550 2.190 ;
        RECT  3.430 0.800 3.540 2.100 ;
        RECT  3.290 0.800 3.430 0.920 ;
        RECT  0.595 1.980 3.430 2.100 ;
        RECT  3.190 1.040 3.310 1.860 ;
        RECT  3.170 0.660 3.290 0.920 ;
        RECT  2.470 1.740 3.190 1.860 ;
        RECT  2.930 0.420 3.050 1.620 ;
        RECT  2.520 0.420 2.930 0.540 ;
        RECT  2.640 1.500 2.930 1.620 ;
        RECT  2.680 0.660 2.800 1.380 ;
        RECT  2.470 1.260 2.680 1.380 ;
        RECT  2.400 0.420 2.520 0.780 ;
        RECT  2.350 1.260 2.470 1.860 ;
        RECT  2.160 0.900 2.420 1.140 ;
        RECT  1.230 0.660 2.400 0.780 ;
        RECT  1.410 1.740 2.350 1.860 ;
        RECT  0.710 0.420 2.180 0.540 ;
        RECT  1.470 0.900 2.160 1.020 ;
        RECT  1.350 0.900 1.470 1.160 ;
        RECT  1.150 1.300 1.410 1.860 ;
        RECT  0.970 1.040 1.350 1.160 ;
        RECT  1.110 0.660 1.230 0.920 ;
        RECT  0.905 0.660 0.970 1.160 ;
        RECT  0.850 0.660 0.905 1.780 ;
        RECT  0.730 1.040 0.850 1.780 ;
        RECT  0.595 0.420 0.710 0.910 ;
        RECT  0.475 0.420 0.595 2.100 ;
    END
END DFFX4AD
MACRO DFFXLAD
    CLASS CORE ;
    FOREIGN DFFXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.950 0.730 6.090 1.700 ;
        RECT  5.895 0.730 5.950 0.900 ;
        RECT  5.930 1.440 5.950 1.700 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 0.730 5.530 1.480 ;
        RECT  5.205 0.730 5.390 0.900 ;
        RECT  5.280 1.340 5.390 1.480 ;
        RECT  5.160 1.340 5.280 1.600 ;
        END
        AntennaDiffArea 0.138 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.740 0.235 1.380 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.705 1.190 1.935 1.610 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.800 -0.210 6.160 0.210 ;
        RECT  5.540 -0.210 5.800 0.435 ;
        RECT  4.635 -0.210 5.540 0.210 ;
        RECT  4.465 -0.210 4.635 0.325 ;
        RECT  3.480 -0.210 4.465 0.210 ;
        RECT  3.220 -0.210 3.480 0.300 ;
        RECT  2.520 -0.210 3.220 0.210 ;
        RECT  2.260 -0.210 2.520 0.300 ;
        RECT  1.790 -0.210 2.260 0.210 ;
        RECT  1.530 -0.210 1.790 0.300 ;
        RECT  0.265 -0.210 1.530 0.210 ;
        RECT  0.095 -0.210 0.265 0.535 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.730 2.310 6.160 2.730 ;
        RECT  5.470 2.020 5.730 2.730 ;
        RECT  4.670 2.310 5.470 2.730 ;
        RECT  4.410 2.060 4.670 2.730 ;
        RECT  3.280 2.310 4.410 2.730 ;
        RECT  3.020 2.220 3.280 2.730 ;
        RECT  2.220 2.310 3.020 2.730 ;
        RECT  1.960 2.220 2.220 2.730 ;
        RECT  1.500 2.310 1.960 2.730 ;
        RECT  1.240 2.220 1.500 2.730 ;
        RECT  0.265 2.310 1.240 2.730 ;
        RECT  0.095 1.595 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.810 1.020 5.830 1.280 ;
        RECT  5.690 1.020 5.810 1.840 ;
        RECT  5.040 1.720 5.690 1.840 ;
        RECT  4.940 0.595 5.040 1.840 ;
        RECT  4.920 0.595 4.940 1.940 ;
        RECT  4.845 0.595 4.920 0.765 ;
        RECT  4.820 1.505 4.920 1.940 ;
        RECT  4.140 1.820 4.820 1.940 ;
        RECT  4.530 0.995 4.790 1.255 ;
        RECT  4.410 0.690 4.530 1.670 ;
        RECT  4.040 0.690 4.410 0.810 ;
        RECT  3.875 1.550 4.410 1.670 ;
        RECT  4.130 0.940 4.260 1.060 ;
        RECT  4.000 0.940 4.130 1.430 ;
        RECT  3.920 0.550 4.040 0.810 ;
        RECT  3.510 1.310 4.000 1.430 ;
        RECT  3.775 0.930 3.880 1.190 ;
        RECT  3.705 1.550 3.875 1.720 ;
        RECT  3.655 0.420 3.775 1.190 ;
        RECT  3.510 1.980 3.770 2.100 ;
        RECT  3.090 0.420 3.655 0.540 ;
        RECT  3.390 0.800 3.510 2.100 ;
        RECT  3.240 0.800 3.390 0.920 ;
        RECT  0.590 1.980 3.390 2.100 ;
        RECT  3.150 1.100 3.270 1.860 ;
        RECT  3.120 0.660 3.240 0.920 ;
        RECT  2.490 1.740 3.150 1.860 ;
        RECT  3.000 0.380 3.090 0.540 ;
        RECT  2.880 0.380 3.000 1.620 ;
        RECT  2.830 0.380 2.880 0.540 ;
        RECT  2.630 1.500 2.880 1.620 ;
        RECT  2.430 0.420 2.830 0.540 ;
        RECT  2.640 0.660 2.760 1.325 ;
        RECT  2.490 1.205 2.640 1.325 ;
        RECT  2.370 1.205 2.490 1.860 ;
        RECT  2.310 0.420 2.430 0.830 ;
        RECT  1.420 1.740 2.370 1.860 ;
        RECT  1.230 0.710 2.310 0.830 ;
        RECT  2.110 0.950 2.230 1.230 ;
        RECT  1.955 0.365 2.125 0.540 ;
        RECT  1.475 0.950 2.110 1.070 ;
        RECT  0.700 0.420 1.955 0.540 ;
        RECT  1.355 0.950 1.475 1.160 ;
        RECT  1.290 1.290 1.420 1.860 ;
        RECT  0.970 1.040 1.355 1.160 ;
        RECT  1.160 1.290 1.290 1.410 ;
        RECT  1.110 0.660 1.230 0.920 ;
        RECT  0.860 0.660 0.970 1.160 ;
        RECT  0.850 0.660 0.860 1.770 ;
        RECT  0.740 1.040 0.850 1.770 ;
        RECT  0.590 0.420 0.700 0.900 ;
        RECT  0.580 0.420 0.590 2.100 ;
        RECT  0.470 0.680 0.580 2.100 ;
    END
END DFFXLAD
MACRO DFFYQX2AD
    CLASS CORE ;
    FOREIGN DFFYQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.930 0.410 6.090 2.015 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.220 1.000 0.340 1.375 ;
        RECT  0.070 1.145 0.220 1.375 ;
        END
        AntennaGateArea 0.146 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.590 1.445 2.160 1.610 ;
        END
        AntennaGateArea 0.133 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 -0.210 6.160 0.210 ;
        RECT  5.545 -0.210 5.715 0.675 ;
        RECT  5.005 -0.210 5.545 0.210 ;
        RECT  4.835 -0.210 5.005 0.420 ;
        RECT  3.780 -0.210 4.835 0.210 ;
        RECT  3.520 -0.210 3.780 0.700 ;
        RECT  2.370 -0.210 3.520 0.210 ;
        RECT  1.850 -0.210 2.370 0.260 ;
        RECT  0.270 -0.210 1.850 0.210 ;
        RECT  0.100 -0.210 0.270 0.785 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 2.310 6.160 2.730 ;
        RECT  5.545 1.845 5.715 2.730 ;
        RECT  4.985 2.310 5.545 2.730 ;
        RECT  4.815 1.945 4.985 2.730 ;
        RECT  3.770 2.310 4.815 2.730 ;
        RECT  3.510 2.210 3.770 2.730 ;
        RECT  2.660 2.310 3.510 2.730 ;
        RECT  2.400 2.210 2.660 2.730 ;
        RECT  1.920 2.310 2.400 2.730 ;
        RECT  1.660 2.010 1.920 2.730 ;
        RECT  0.270 2.310 1.660 2.730 ;
        RECT  0.100 1.600 0.270 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.680 0.820 5.800 1.695 ;
        RECT  5.365 0.820 5.680 0.940 ;
        RECT  4.790 1.525 5.680 1.695 ;
        RECT  5.030 1.065 5.535 1.235 ;
        RECT  5.195 0.735 5.365 0.940 ;
        RECT  4.910 0.620 5.030 1.235 ;
        RECT  4.330 0.620 4.910 0.740 ;
        RECT  4.670 1.120 4.790 1.695 ;
        RECT  4.330 1.970 4.590 2.190 ;
        RECT  4.290 0.330 4.550 0.500 ;
        RECT  4.210 0.620 4.330 1.730 ;
        RECT  4.040 1.970 4.330 2.090 ;
        RECT  4.020 0.380 4.290 0.500 ;
        RECT  4.140 0.620 4.210 0.740 ;
        RECT  4.020 0.820 4.040 2.090 ;
        RECT  3.920 0.380 4.020 2.090 ;
        RECT  3.900 0.380 3.920 0.940 ;
        RECT  2.235 1.970 3.920 2.090 ;
        RECT  3.560 0.820 3.900 0.940 ;
        RECT  3.680 1.060 3.800 1.850 ;
        RECT  2.970 1.730 3.680 1.850 ;
        RECT  3.440 0.820 3.560 1.320 ;
        RECT  3.350 1.060 3.440 1.320 ;
        RECT  3.210 1.490 3.390 1.610 ;
        RECT  3.270 0.640 3.320 0.900 ;
        RECT  3.210 0.330 3.270 0.900 ;
        RECT  3.090 0.330 3.210 1.610 ;
        RECT  3.010 0.330 3.090 0.610 ;
        RECT  2.750 0.490 3.010 0.610 ;
        RECT  2.850 0.730 2.970 1.850 ;
        RECT  2.780 1.505 2.850 1.850 ;
        RECT  2.400 1.505 2.780 1.625 ;
        RECT  2.630 0.380 2.750 0.610 ;
        RECT  2.610 0.890 2.730 1.280 ;
        RECT  1.495 0.380 2.630 0.500 ;
        RECT  1.175 0.890 2.610 1.010 ;
        RECT  1.205 0.650 2.400 0.770 ;
        RECT  2.280 1.200 2.400 1.625 ;
        RECT  1.540 1.200 2.280 1.320 ;
        RECT  2.065 1.770 2.235 2.090 ;
        RECT  1.075 1.770 2.065 1.890 ;
        RECT  1.325 0.330 1.495 0.500 ;
        RECT  1.175 1.480 1.265 1.650 ;
        RECT  1.085 0.380 1.205 0.770 ;
        RECT  1.005 0.890 1.175 1.650 ;
        RECT  0.585 0.380 1.085 0.500 ;
        RECT  0.905 1.770 1.075 2.190 ;
        RECT  0.965 0.890 1.005 1.010 ;
        RECT  0.835 1.480 1.005 1.650 ;
        RECT  0.845 0.650 0.965 1.010 ;
        RECT  0.715 1.770 0.905 1.890 ;
        RECT  0.705 0.650 0.845 0.770 ;
        RECT  0.715 0.890 0.725 1.150 ;
        RECT  0.595 0.890 0.715 1.890 ;
        RECT  0.585 0.890 0.595 1.150 ;
        RECT  0.465 0.380 0.585 1.150 ;
    END
END DFFYQX2AD
MACRO DLY1X1AD
    CLASS CORE ;
    FOREIGN DLY1X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.650 2.450 1.905 ;
        RECT  2.280 0.650 2.310 0.910 ;
        RECT  2.280 1.385 2.310 1.905 ;
        END
        AntennaDiffArea 0.2 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.515 1.390 ;
        RECT  0.325 1.095 0.350 1.390 ;
        END
        AntennaGateArea 0.0594 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 -0.210 2.520 0.210 ;
        RECT  1.955 -0.210 2.125 0.325 ;
        RECT  0.635 -0.210 1.955 0.210 ;
        RECT  0.465 -0.210 0.635 0.380 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 2.310 2.520 2.730 ;
        RECT  1.955 2.195 2.125 2.730 ;
        RECT  0.635 2.310 1.955 2.730 ;
        RECT  0.465 1.975 0.635 2.730 ;
        RECT  0.000 2.310 0.465 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.065 1.010 2.190 1.270 ;
        RECT  1.895 0.445 2.065 2.075 ;
        RECT  1.460 0.445 1.895 0.615 ;
        RECT  1.265 1.905 1.895 2.075 ;
        RECT  1.630 0.750 1.750 1.530 ;
        RECT  1.280 1.055 1.630 1.225 ;
        RECT  1.200 0.330 1.460 0.615 ;
        RECT  1.245 0.800 1.280 1.225 ;
        RECT  1.075 0.800 1.245 1.630 ;
        RECT  0.890 1.150 0.915 1.700 ;
        RECT  0.770 1.080 0.890 1.700 ;
        RECT  0.745 1.150 0.770 1.700 ;
        RECT  0.205 1.530 0.745 1.700 ;
        RECT  0.205 0.630 0.230 0.890 ;
        RECT  0.085 0.630 0.205 1.700 ;
    END
END DLY1X1AD
MACRO DLY1X4AD
    CLASS CORE ;
    FOREIGN DLY1X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.705 0.440 2.730 1.235 ;
        RECT  2.555 0.440 2.705 2.075 ;
        RECT  2.495 0.440 2.555 0.870 ;
        RECT  2.465 1.645 2.555 2.075 ;
        END
        AntennaDiffArea 0.391 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.535 1.375 ;
        RECT  0.325 0.975 0.350 1.375 ;
        END
        AntennaGateArea 0.1004 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.305 -0.210 3.080 0.210 ;
        RECT  2.135 -0.210 2.305 0.525 ;
        RECT  0.635 -0.210 2.135 0.210 ;
        RECT  0.465 -0.210 0.635 0.255 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.995 2.310 3.080 2.730 ;
        RECT  2.825 1.645 2.995 2.730 ;
        RECT  2.205 2.310 2.825 2.730 ;
        RECT  2.035 2.165 2.205 2.730 ;
        RECT  0.635 2.310 2.035 2.730 ;
        RECT  0.465 2.195 0.635 2.730 ;
        RECT  0.000 2.310 0.465 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  2.190 0.675 2.360 1.580 ;
        RECT  1.435 0.675 2.190 0.845 ;
        RECT  1.605 1.410 2.190 1.580 ;
        RECT  1.265 1.055 1.935 1.225 ;
        RECT  1.435 1.410 1.605 1.840 ;
        RECT  1.095 0.645 1.265 1.905 ;
        RECT  0.765 1.055 0.935 1.665 ;
        RECT  0.255 1.495 0.765 1.665 ;
        RECT  0.205 1.495 0.255 1.925 ;
        RECT  0.205 0.605 0.230 0.865 ;
        RECT  0.085 0.605 0.205 1.925 ;
    END
END DLY1X4AD
MACRO DLY2X1AD
    CLASS CORE ;
    FOREIGN DLY2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.650 2.450 1.905 ;
        RECT  2.280 0.650 2.310 0.910 ;
        RECT  2.280 1.385 2.310 1.905 ;
        END
        AntennaDiffArea 0.2 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.515 1.390 ;
        RECT  0.325 1.095 0.350 1.390 ;
        END
        AntennaGateArea 0.0594 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 -0.210 2.520 0.210 ;
        RECT  1.955 -0.210 2.125 0.325 ;
        RECT  0.635 -0.210 1.955 0.210 ;
        RECT  0.465 -0.210 0.635 0.380 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 2.310 2.520 2.730 ;
        RECT  1.955 2.195 2.125 2.730 ;
        RECT  0.635 2.310 1.955 2.730 ;
        RECT  0.465 1.975 0.635 2.730 ;
        RECT  0.000 2.310 0.465 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.065 1.010 2.190 1.270 ;
        RECT  1.895 0.445 2.065 2.075 ;
        RECT  1.460 0.445 1.895 0.615 ;
        RECT  1.265 1.905 1.895 2.075 ;
        RECT  1.630 0.750 1.750 1.530 ;
        RECT  1.280 1.055 1.630 1.225 ;
        RECT  1.200 0.330 1.460 0.615 ;
        RECT  1.245 0.800 1.280 1.225 ;
        RECT  1.075 0.800 1.245 1.630 ;
        RECT  0.890 1.150 0.915 1.700 ;
        RECT  0.770 1.080 0.890 1.700 ;
        RECT  0.745 1.150 0.770 1.700 ;
        RECT  0.205 1.530 0.745 1.700 ;
        RECT  0.205 0.630 0.230 0.890 ;
        RECT  0.085 0.630 0.205 1.700 ;
    END
END DLY2X1AD
MACRO DLY2X4AD
    CLASS CORE ;
    FOREIGN DLY2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.705 0.440 2.730 1.235 ;
        RECT  2.555 0.440 2.705 2.075 ;
        RECT  2.495 0.440 2.555 0.870 ;
        RECT  2.465 1.645 2.555 2.075 ;
        END
        AntennaDiffArea 0.391 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.535 1.375 ;
        RECT  0.325 0.975 0.350 1.375 ;
        END
        AntennaGateArea 0.1004 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.305 -0.210 3.080 0.210 ;
        RECT  2.135 -0.210 2.305 0.525 ;
        RECT  0.635 -0.210 2.135 0.210 ;
        RECT  0.465 -0.210 0.635 0.255 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.995 2.310 3.080 2.730 ;
        RECT  2.825 1.645 2.995 2.730 ;
        RECT  2.205 2.310 2.825 2.730 ;
        RECT  2.035 2.165 2.205 2.730 ;
        RECT  0.635 2.310 2.035 2.730 ;
        RECT  0.465 2.195 0.635 2.730 ;
        RECT  0.000 2.310 0.465 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  2.190 0.675 2.360 1.580 ;
        RECT  1.435 0.675 2.190 0.845 ;
        RECT  1.605 1.410 2.190 1.580 ;
        RECT  1.265 1.055 1.935 1.225 ;
        RECT  1.435 1.410 1.605 1.840 ;
        RECT  1.095 0.645 1.265 1.905 ;
        RECT  0.765 1.055 0.935 1.665 ;
        RECT  0.255 1.495 0.765 1.665 ;
        RECT  0.205 1.495 0.255 1.925 ;
        RECT  0.205 0.605 0.230 0.865 ;
        RECT  0.085 0.605 0.205 1.925 ;
    END
END DLY2X4AD
MACRO DLY3X1AD
    CLASS CORE ;
    FOREIGN DLY3X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.650 2.450 1.905 ;
        RECT  2.280 0.650 2.310 0.910 ;
        RECT  2.280 1.385 2.310 1.905 ;
        END
        AntennaDiffArea 0.2 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.515 1.390 ;
        RECT  0.325 1.095 0.350 1.390 ;
        END
        AntennaGateArea 0.0594 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 -0.210 2.520 0.210 ;
        RECT  1.955 -0.210 2.125 0.325 ;
        RECT  0.635 -0.210 1.955 0.210 ;
        RECT  0.465 -0.210 0.635 0.380 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 2.310 2.520 2.730 ;
        RECT  1.955 2.195 2.125 2.730 ;
        RECT  0.635 2.310 1.955 2.730 ;
        RECT  0.465 1.975 0.635 2.730 ;
        RECT  0.000 2.310 0.465 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.065 1.010 2.190 1.270 ;
        RECT  1.895 0.445 2.065 2.075 ;
        RECT  1.460 0.445 1.895 0.615 ;
        RECT  1.265 1.905 1.895 2.075 ;
        RECT  1.630 0.750 1.750 1.530 ;
        RECT  1.280 1.055 1.630 1.225 ;
        RECT  1.200 0.330 1.460 0.615 ;
        RECT  1.245 0.800 1.280 1.225 ;
        RECT  1.075 0.800 1.245 1.630 ;
        RECT  0.890 1.150 0.915 1.700 ;
        RECT  0.770 1.080 0.890 1.700 ;
        RECT  0.745 1.150 0.770 1.700 ;
        RECT  0.205 1.530 0.745 1.700 ;
        RECT  0.205 0.630 0.230 0.890 ;
        RECT  0.085 0.630 0.205 1.700 ;
    END
END DLY3X1AD
MACRO DLY3X4AD
    CLASS CORE ;
    FOREIGN DLY3X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.705 0.440 2.730 1.235 ;
        RECT  2.555 0.440 2.705 2.075 ;
        RECT  2.495 0.440 2.555 0.870 ;
        RECT  2.465 1.645 2.555 2.075 ;
        END
        AntennaDiffArea 0.391 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.535 1.375 ;
        RECT  0.325 0.975 0.350 1.375 ;
        END
        AntennaGateArea 0.1004 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.305 -0.210 3.080 0.210 ;
        RECT  2.135 -0.210 2.305 0.525 ;
        RECT  0.635 -0.210 2.135 0.210 ;
        RECT  0.465 -0.210 0.635 0.255 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.995 2.310 3.080 2.730 ;
        RECT  2.825 1.645 2.995 2.730 ;
        RECT  2.205 2.310 2.825 2.730 ;
        RECT  2.035 2.165 2.205 2.730 ;
        RECT  0.635 2.310 2.035 2.730 ;
        RECT  0.465 2.195 0.635 2.730 ;
        RECT  0.000 2.310 0.465 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  2.190 0.675 2.360 1.580 ;
        RECT  1.435 0.675 2.190 0.845 ;
        RECT  1.605 1.410 2.190 1.580 ;
        RECT  1.265 1.055 1.935 1.225 ;
        RECT  1.435 1.410 1.605 1.840 ;
        RECT  1.095 0.645 1.265 1.905 ;
        RECT  0.765 1.055 0.935 1.665 ;
        RECT  0.255 1.495 0.765 1.665 ;
        RECT  0.205 1.495 0.255 1.925 ;
        RECT  0.205 0.605 0.230 0.865 ;
        RECT  0.085 0.605 0.205 1.925 ;
    END
END DLY3X4AD
MACRO DLY4X1AD
    CLASS CORE ;
    FOREIGN DLY4X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.650 2.450 1.905 ;
        RECT  2.280 0.650 2.310 0.910 ;
        RECT  2.280 1.385 2.310 1.905 ;
        END
        AntennaDiffArea 0.2 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.515 1.390 ;
        RECT  0.325 1.095 0.350 1.390 ;
        END
        AntennaGateArea 0.0594 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 -0.210 2.520 0.210 ;
        RECT  1.955 -0.210 2.125 0.325 ;
        RECT  0.635 -0.210 1.955 0.210 ;
        RECT  0.465 -0.210 0.635 0.380 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 2.310 2.520 2.730 ;
        RECT  1.955 2.195 2.125 2.730 ;
        RECT  0.635 2.310 1.955 2.730 ;
        RECT  0.465 1.975 0.635 2.730 ;
        RECT  0.000 2.310 0.465 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.065 1.010 2.190 1.270 ;
        RECT  1.895 0.445 2.065 2.075 ;
        RECT  1.460 0.445 1.895 0.615 ;
        RECT  1.265 1.905 1.895 2.075 ;
        RECT  1.630 0.750 1.750 1.530 ;
        RECT  1.280 1.055 1.630 1.225 ;
        RECT  1.200 0.330 1.460 0.615 ;
        RECT  1.245 0.800 1.280 1.225 ;
        RECT  1.075 0.800 1.245 1.630 ;
        RECT  0.890 1.150 0.915 1.700 ;
        RECT  0.770 1.080 0.890 1.700 ;
        RECT  0.745 1.150 0.770 1.700 ;
        RECT  0.205 1.530 0.745 1.700 ;
        RECT  0.205 0.630 0.230 0.890 ;
        RECT  0.085 0.630 0.205 1.700 ;
    END
END DLY4X1AD
MACRO DLY4X4AD
    CLASS CORE ;
    FOREIGN DLY4X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.705 0.440 2.730 1.235 ;
        RECT  2.555 0.440 2.705 2.075 ;
        RECT  2.495 0.440 2.555 0.870 ;
        RECT  2.465 1.645 2.555 2.075 ;
        END
        AntennaDiffArea 0.391 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.535 1.375 ;
        RECT  0.325 0.975 0.350 1.375 ;
        END
        AntennaGateArea 0.1004 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.305 -0.210 3.080 0.210 ;
        RECT  2.135 -0.210 2.305 0.525 ;
        RECT  0.635 -0.210 2.135 0.210 ;
        RECT  0.465 -0.210 0.635 0.255 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.995 2.310 3.080 2.730 ;
        RECT  2.825 1.645 2.995 2.730 ;
        RECT  2.205 2.310 2.825 2.730 ;
        RECT  2.035 2.165 2.205 2.730 ;
        RECT  0.635 2.310 2.035 2.730 ;
        RECT  0.465 2.195 0.635 2.730 ;
        RECT  0.000 2.310 0.465 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  2.190 0.675 2.360 1.580 ;
        RECT  1.435 0.675 2.190 0.845 ;
        RECT  1.605 1.410 2.190 1.580 ;
        RECT  1.265 1.055 1.935 1.225 ;
        RECT  1.435 1.410 1.605 1.840 ;
        RECT  1.095 0.645 1.265 1.905 ;
        RECT  0.765 1.055 0.935 1.665 ;
        RECT  0.255 1.495 0.765 1.665 ;
        RECT  0.205 1.495 0.255 1.925 ;
        RECT  0.205 0.605 0.230 0.865 ;
        RECT  0.085 0.605 0.205 1.925 ;
    END
END DLY4X4AD
MACRO EDFFHQX1AD
    CLASS CORE ;
    FOREIGN EDFFHQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.560 1.145 8.610 1.375 ;
        RECT  8.440 0.645 8.560 1.860 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.740 1.375 3.910 1.495 ;
        RECT  3.620 1.040 3.740 1.495 ;
        RECT  3.260 1.040 3.620 1.160 ;
        RECT  3.140 0.900 3.260 1.620 ;
        RECT  3.090 0.900 3.140 1.160 ;
        RECT  1.890 1.500 3.140 1.620 ;
        RECT  1.770 1.145 1.890 1.620 ;
        RECT  1.600 1.145 1.770 1.445 ;
        END
        AntennaGateArea 0.101 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.495 0.860 2.730 1.120 ;
        END
        AntennaGateArea 0.095 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.025 0.570 1.375 ;
        END
        AntennaGateArea 0.131 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.225 -0.210 8.680 0.210 ;
        RECT  8.055 -0.210 8.225 0.900 ;
        RECT  7.570 -0.210 8.055 0.210 ;
        RECT  7.450 -0.210 7.570 0.610 ;
        RECT  6.090 -0.210 7.450 0.210 ;
        RECT  5.830 -0.210 6.090 0.260 ;
        RECT  4.320 -0.210 5.830 0.210 ;
        RECT  3.800 -0.210 4.320 0.260 ;
        RECT  2.395 -0.210 3.800 0.210 ;
        RECT  2.275 -0.210 2.395 0.370 ;
        RECT  1.100 -0.210 2.275 0.210 ;
        RECT  0.580 -0.210 1.100 0.300 ;
        RECT  0.000 -0.210 0.580 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.195 2.310 8.680 2.730 ;
        RECT  7.675 2.220 8.195 2.730 ;
        RECT  5.620 2.310 7.675 2.730 ;
        RECT  5.360 2.220 5.620 2.730 ;
        RECT  4.480 2.310 5.360 2.730 ;
        RECT  4.220 2.220 4.480 2.730 ;
        RECT  2.700 2.310 4.220 2.730 ;
        RECT  2.440 2.220 2.700 2.730 ;
        RECT  2.050 2.310 2.440 2.730 ;
        RECT  1.790 2.220 2.050 2.730 ;
        RECT  0.610 2.310 1.790 2.730 ;
        RECT  0.350 1.975 0.610 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.680 2.520 ;
        LAYER M1 ;
        RECT  8.155 1.020 8.275 2.090 ;
        RECT  7.895 1.020 8.155 1.280 ;
        RECT  7.160 1.970 8.155 2.090 ;
        RECT  7.770 0.755 7.910 0.875 ;
        RECT  7.770 1.430 7.910 1.550 ;
        RECT  7.650 0.755 7.770 1.550 ;
        RECT  7.640 1.330 7.650 1.550 ;
        RECT  7.090 1.330 7.640 1.450 ;
        RECT  7.210 0.380 7.330 1.160 ;
        RECT  6.670 0.380 7.210 0.500 ;
        RECT  7.040 1.590 7.160 2.150 ;
        RECT  6.970 0.620 7.090 1.450 ;
        RECT  6.775 1.590 7.040 1.710 ;
        RECT  4.220 0.620 6.970 0.740 ;
        RECT  6.100 1.830 6.870 1.950 ;
        RECT  6.775 0.875 6.825 1.045 ;
        RECT  6.655 0.875 6.775 1.710 ;
        RECT  6.410 0.330 6.670 0.500 ;
        RECT  6.220 1.590 6.655 1.710 ;
        RECT  6.100 0.900 6.490 1.020 ;
        RECT  5.550 0.380 6.410 0.500 ;
        RECT  5.860 2.070 6.250 2.190 ;
        RECT  5.980 0.900 6.100 1.950 ;
        RECT  5.650 0.900 5.980 1.030 ;
        RECT  4.500 1.740 5.980 1.860 ;
        RECT  5.740 1.980 5.860 2.190 ;
        RECT  5.690 1.150 5.810 1.410 ;
        RECT  4.930 1.980 5.740 2.100 ;
        RECT  5.410 1.220 5.690 1.340 ;
        RECT  5.290 0.330 5.550 0.500 ;
        RECT  5.290 0.860 5.410 1.620 ;
        RECT  2.635 0.380 5.290 0.500 ;
        RECT  5.060 0.860 5.290 0.980 ;
        RECT  4.820 1.500 5.290 1.620 ;
        RECT  4.865 1.200 5.170 1.320 ;
        RECT  4.670 1.980 4.930 2.190 ;
        RECT  4.745 1.110 4.865 1.320 ;
        RECT  4.180 1.110 4.745 1.230 ;
        RECT  3.980 1.980 4.670 2.100 ;
        RECT  4.380 1.350 4.500 1.860 ;
        RECT  4.100 0.620 4.220 0.990 ;
        RECT  4.060 1.110 4.180 1.760 ;
        RECT  3.980 1.110 4.060 1.230 ;
        RECT  3.740 1.640 4.060 1.760 ;
        RECT  3.860 0.620 3.980 1.230 ;
        RECT  3.860 1.980 3.980 2.140 ;
        RECT  3.140 0.620 3.860 0.740 ;
        RECT  3.500 2.020 3.860 2.140 ;
        RECT  3.620 1.640 3.740 1.900 ;
        RECT  3.380 1.280 3.500 1.860 ;
        RECT  3.380 1.980 3.500 2.140 ;
        RECT  1.590 1.740 3.380 1.860 ;
        RECT  1.250 1.980 3.380 2.100 ;
        RECT  2.970 0.620 3.020 0.740 ;
        RECT  2.970 1.260 3.020 1.380 ;
        RECT  2.850 0.620 2.970 1.380 ;
        RECT  2.760 0.620 2.850 0.740 ;
        RECT  2.760 1.260 2.850 1.380 ;
        RECT  2.515 0.380 2.635 0.710 ;
        RECT  2.170 0.590 2.515 0.710 ;
        RECT  2.170 1.260 2.310 1.380 ;
        RECT  2.050 0.590 2.170 1.380 ;
        RECT  1.825 0.590 2.050 0.780 ;
        RECT  1.170 0.660 1.825 0.780 ;
        RECT  1.400 0.350 1.800 0.470 ;
        RECT  1.410 0.900 1.660 1.020 ;
        RECT  1.470 1.575 1.590 1.860 ;
        RECT  1.410 1.575 1.470 1.695 ;
        RECT  1.290 0.900 1.410 1.695 ;
        RECT  1.280 0.350 1.400 0.540 ;
        RECT  0.240 0.420 1.280 0.540 ;
        RECT  1.110 1.815 1.250 2.100 ;
        RECT  1.050 0.660 1.170 1.330 ;
        RECT  0.990 1.450 1.110 2.100 ;
        RECT  0.990 1.070 1.050 1.330 ;
        RECT  0.870 1.450 0.990 1.570 ;
        RECT  0.870 0.690 0.930 0.950 ;
        RECT  0.810 0.690 0.870 1.570 ;
        RECT  0.750 0.830 0.810 1.570 ;
        RECT  0.215 0.420 0.240 0.950 ;
        RECT  0.215 1.440 0.240 1.700 ;
        RECT  0.120 0.420 0.215 1.700 ;
        RECT  0.095 0.735 0.120 1.700 ;
    END
END EDFFHQX1AD
MACRO EDFFHQX2AD
    CLASS CORE ;
    FOREIGN EDFFHQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.850 1.145 8.890 1.375 ;
        RECT  8.730 0.370 8.850 2.155 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 1.440 3.875 1.560 ;
        RECT  3.430 0.865 3.590 1.095 ;
        RECT  3.310 0.865 3.430 1.620 ;
        RECT  3.150 0.865 3.310 1.095 ;
        RECT  1.855 1.500 3.310 1.620 ;
        RECT  1.735 1.150 1.855 1.620 ;
        RECT  1.535 1.150 1.735 1.410 ;
        END
        AntennaGateArea 0.112 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.300 0.860 2.685 1.120 ;
        END
        AntennaGateArea 0.14 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.060 0.805 1.445 ;
        END
        AntennaGateArea 0.143 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.515 -0.210 8.960 0.210 ;
        RECT  8.255 -0.210 8.515 0.450 ;
        RECT  7.830 -0.210 8.255 0.210 ;
        RECT  7.670 -0.210 7.830 0.690 ;
        RECT  5.990 -0.210 7.670 0.210 ;
        RECT  5.730 -0.210 5.990 0.260 ;
        RECT  4.345 -0.210 5.730 0.210 ;
        RECT  4.225 -0.210 4.345 0.370 ;
        RECT  2.425 -0.210 4.225 0.210 ;
        RECT  2.305 -0.210 2.425 0.370 ;
        RECT  1.100 -0.210 2.305 0.210 ;
        RECT  0.580 -0.210 1.100 0.300 ;
        RECT  0.000 -0.210 0.580 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.530 2.310 8.960 2.730 ;
        RECT  8.010 2.020 8.530 2.730 ;
        RECT  6.430 2.310 8.010 2.730 ;
        RECT  6.170 2.220 6.430 2.730 ;
        RECT  5.670 2.310 6.170 2.730 ;
        RECT  5.410 2.220 5.670 2.730 ;
        RECT  4.415 2.310 5.410 2.730 ;
        RECT  4.155 2.255 4.415 2.730 ;
        RECT  2.555 2.310 4.155 2.730 ;
        RECT  2.295 2.290 2.555 2.730 ;
        RECT  1.955 2.310 2.295 2.730 ;
        RECT  1.695 2.220 1.955 2.730 ;
        RECT  0.635 2.310 1.695 2.730 ;
        RECT  0.375 1.930 0.635 2.730 ;
        RECT  0.000 2.310 0.375 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.960 2.520 ;
        LAYER M1 ;
        RECT  8.470 1.050 8.610 1.170 ;
        RECT  8.350 1.050 8.470 1.850 ;
        RECT  7.555 1.730 8.350 1.850 ;
        RECT  8.060 0.690 8.180 1.610 ;
        RECT  7.870 1.050 8.060 1.380 ;
        RECT  7.310 1.260 7.870 1.380 ;
        RECT  7.550 1.020 7.720 1.140 ;
        RECT  7.505 1.730 7.555 2.045 ;
        RECT  7.430 0.380 7.550 1.140 ;
        RECT  7.385 1.500 7.505 2.045 ;
        RECT  7.005 0.380 7.430 0.500 ;
        RECT  7.070 1.500 7.385 1.620 ;
        RECT  7.190 0.620 7.310 1.380 ;
        RECT  6.320 1.740 7.240 1.860 ;
        RECT  4.830 0.620 7.190 0.740 ;
        RECT  6.950 0.860 7.070 1.620 ;
        RECT  6.745 0.330 7.005 0.500 ;
        RECT  6.550 0.860 6.950 0.980 ;
        RECT  6.620 1.500 6.950 1.620 ;
        RECT  5.410 0.380 6.745 0.500 ;
        RECT  4.850 1.980 6.690 2.100 ;
        RECT  6.320 0.900 6.390 1.020 ;
        RECT  6.200 0.900 6.320 1.860 ;
        RECT  5.750 0.900 6.200 1.020 ;
        RECT  4.460 1.740 6.200 1.860 ;
        RECT  5.340 1.310 6.045 1.430 ;
        RECT  5.490 0.900 5.750 1.055 ;
        RECT  5.150 0.330 5.410 0.500 ;
        RECT  5.220 0.900 5.340 1.620 ;
        RECT  4.960 0.860 5.220 1.020 ;
        RECT  4.780 1.500 5.220 1.620 ;
        RECT  4.585 0.380 5.150 0.500 ;
        RECT  5.055 1.200 5.100 1.320 ;
        RECT  4.840 1.140 5.055 1.320 ;
        RECT  4.590 1.980 4.850 2.190 ;
        RECT  4.155 1.140 4.840 1.260 ;
        RECT  4.710 0.620 4.830 1.020 ;
        RECT  4.000 0.900 4.710 1.020 ;
        RECT  1.155 1.980 4.590 2.100 ;
        RECT  4.465 0.380 4.585 0.765 ;
        RECT  4.105 0.645 4.465 0.765 ;
        RECT  4.340 1.380 4.460 1.860 ;
        RECT  4.275 1.380 4.340 1.550 ;
        RECT  4.035 1.140 4.155 1.850 ;
        RECT  3.985 0.380 4.105 0.765 ;
        RECT  3.865 1.140 4.035 1.260 ;
        RECT  3.495 1.730 4.035 1.850 ;
        RECT  2.665 0.380 3.985 0.500 ;
        RECT  3.745 0.620 3.865 1.260 ;
        RECT  3.235 0.620 3.745 0.740 ;
        RECT  3.030 1.260 3.190 1.380 ;
        RECT  1.575 1.740 3.135 1.860 ;
        RECT  3.030 0.620 3.070 0.740 ;
        RECT  2.910 0.620 3.030 1.380 ;
        RECT  2.810 0.620 2.910 0.740 ;
        RECT  2.545 0.380 2.665 0.640 ;
        RECT  2.125 0.520 2.545 0.640 ;
        RECT  2.125 1.260 2.265 1.380 ;
        RECT  2.005 0.520 2.125 1.380 ;
        RECT  1.925 0.520 2.005 0.780 ;
        RECT  1.175 0.660 1.925 0.780 ;
        RECT  0.230 0.420 1.805 0.540 ;
        RECT  1.415 0.900 1.625 1.020 ;
        RECT  1.455 1.610 1.575 1.860 ;
        RECT  1.415 1.610 1.455 1.730 ;
        RECT  1.295 0.900 1.415 1.730 ;
        RECT  1.055 0.660 1.175 1.455 ;
        RECT  1.035 1.605 1.155 2.100 ;
        RECT  0.965 1.195 1.055 1.455 ;
        RECT  0.510 1.605 1.035 1.725 ;
        RECT  0.780 0.680 0.900 0.940 ;
        RECT  0.510 0.820 0.780 0.940 ;
        RECT  0.390 0.820 0.510 1.725 ;
        RECT  0.110 0.420 0.230 1.755 ;
    END
END EDFFHQX2AD
MACRO EDFFHQX4AD
    CLASS CORE ;
    FOREIGN EDFFHQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.315 1.005 11.505 1.515 ;
        RECT  11.145 0.385 11.315 2.120 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.945 1.125 2.065 1.890 ;
        RECT  1.705 1.710 1.945 1.890 ;
        RECT  0.830 1.710 1.705 1.830 ;
        RECT  0.710 1.710 0.830 2.135 ;
        RECT  0.385 2.000 0.710 2.135 ;
        RECT  0.125 2.000 0.385 2.175 ;
        END
        AntennaGateArea 0.152 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.820 1.055 1.030 1.225 ;
        RECT  0.570 0.910 0.820 1.225 ;
        END
        AntennaGateArea 0.225 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.105 0.910 3.425 1.180 ;
        END
        AntennaGateArea 0.204 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.675 -0.210 11.760 0.210 ;
        RECT  11.505 -0.210 11.675 0.840 ;
        RECT  11.000 -0.210 11.505 0.210 ;
        RECT  10.740 -0.210 11.000 0.500 ;
        RECT  10.025 -0.210 10.740 0.210 ;
        RECT  9.505 -0.210 10.025 0.500 ;
        RECT  7.465 -0.210 9.505 0.210 ;
        RECT  7.205 -0.210 7.465 0.260 ;
        RECT  6.120 -0.210 7.205 0.210 ;
        RECT  5.600 -0.210 6.120 0.260 ;
        RECT  4.770 -0.210 5.600 0.210 ;
        RECT  4.250 -0.210 4.770 0.260 ;
        RECT  3.360 -0.210 4.250 0.210 ;
        RECT  3.100 -0.210 3.360 0.260 ;
        RECT  2.740 -0.210 3.100 0.210 ;
        RECT  2.480 -0.210 2.740 0.260 ;
        RECT  0.885 -0.210 2.480 0.210 ;
        RECT  0.365 -0.210 0.885 0.330 ;
        RECT  0.000 -0.210 0.365 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.675 2.310 11.760 2.730 ;
        RECT  11.505 1.680 11.675 2.730 ;
        RECT  10.955 2.310 11.505 2.730 ;
        RECT  10.785 1.950 10.955 2.730 ;
        RECT  10.430 2.310 10.785 2.730 ;
        RECT  10.260 1.950 10.430 2.730 ;
        RECT  7.840 2.310 10.260 2.730 ;
        RECT  7.580 2.260 7.840 2.730 ;
        RECT  7.060 2.310 7.580 2.730 ;
        RECT  6.800 2.260 7.060 2.730 ;
        RECT  4.755 2.310 6.800 2.730 ;
        RECT  4.235 2.260 4.755 2.730 ;
        RECT  2.660 2.310 4.235 2.730 ;
        RECT  2.490 1.995 2.660 2.730 ;
        RECT  1.260 2.310 2.490 2.730 ;
        RECT  1.255 1.995 1.260 2.730 ;
        RECT  0.995 1.970 1.255 2.730 ;
        RECT  0.680 2.310 0.995 2.730 ;
        RECT  0.420 2.290 0.680 2.730 ;
        RECT  0.000 2.310 0.420 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.760 2.520 ;
        LAYER M1 ;
        RECT  10.905 0.620 11.025 1.600 ;
        RECT  10.335 0.620 10.905 0.880 ;
        RECT  10.595 1.430 10.905 1.600 ;
        RECT  10.135 1.050 10.785 1.220 ;
        RECT  10.475 1.430 10.595 1.780 ;
        RECT  10.140 1.660 10.475 1.780 ;
        RECT  9.265 0.620 10.335 0.740 ;
        RECT  9.880 1.660 10.140 2.020 ;
        RECT  10.015 0.860 10.135 1.540 ;
        RECT  8.935 0.860 10.015 0.980 ;
        RECT  8.835 1.420 10.015 1.540 ;
        RECT  8.110 1.140 9.895 1.260 ;
        RECT  6.075 2.020 9.670 2.140 ;
        RECT  7.800 1.745 9.455 1.865 ;
        RECT  9.145 0.380 9.265 0.740 ;
        RECT  2.545 0.380 9.145 0.500 ;
        RECT  8.810 0.620 8.935 0.980 ;
        RECT  8.340 0.620 8.810 0.740 ;
        RECT  7.990 0.660 8.110 1.260 ;
        RECT  4.610 0.660 7.990 0.780 ;
        RECT  7.630 0.955 7.800 1.865 ;
        RECT  6.820 1.745 7.630 1.865 ;
        RECT  7.230 1.000 7.350 1.510 ;
        RECT  6.580 1.000 7.230 1.120 ;
        RECT  7.080 1.390 7.230 1.510 ;
        RECT  6.700 1.305 6.820 1.865 ;
        RECT  6.460 1.000 6.580 1.550 ;
        RECT  6.365 1.430 6.460 1.550 ;
        RECT  6.195 1.430 6.365 1.840 ;
        RECT  5.360 1.430 6.195 1.550 ;
        RECT  5.955 1.685 6.075 2.140 ;
        RECT  5.110 0.965 5.970 1.085 ;
        RECT  5.110 1.685 5.955 1.805 ;
        RECT  5.655 1.930 5.775 2.190 ;
        RECT  2.900 2.020 5.655 2.140 ;
        RECT  4.990 0.965 5.110 1.805 ;
        RECT  4.370 1.685 4.990 1.805 ;
        RECT  4.490 0.660 4.610 1.520 ;
        RECT  3.870 0.660 4.490 0.780 ;
        RECT  4.130 1.400 4.490 1.520 ;
        RECT  4.250 1.685 4.370 1.900 ;
        RECT  3.890 0.965 4.325 1.135 ;
        RECT  3.140 1.780 4.250 1.900 ;
        RECT  4.010 1.400 4.130 1.660 ;
        RECT  3.510 1.540 4.010 1.660 ;
        RECT  3.750 0.965 3.890 1.420 ;
        RECT  3.630 0.625 3.750 1.420 ;
        RECT  3.490 0.625 3.630 0.745 ;
        RECT  3.390 1.400 3.510 1.660 ;
        RECT  3.020 1.495 3.140 1.900 ;
        RECT  2.905 0.640 3.120 0.760 ;
        RECT  2.905 1.495 3.020 1.615 ;
        RECT  2.785 0.640 2.905 1.615 ;
        RECT  2.780 1.735 2.900 2.140 ;
        RECT  2.305 1.735 2.780 1.855 ;
        RECT  2.425 0.380 2.545 1.190 ;
        RECT  2.185 0.760 2.305 2.145 ;
        RECT  2.050 0.760 2.185 0.880 ;
        RECT  1.835 2.025 2.185 2.145 ;
        RECT  1.880 0.635 2.050 0.880 ;
        RECT  1.735 0.330 1.905 0.450 ;
        RECT  1.615 0.330 1.735 1.330 ;
        RECT  0.255 0.470 1.615 0.590 ;
        RECT  1.475 1.170 1.615 1.330 ;
        RECT  1.320 1.470 1.615 1.590 ;
        RECT  1.200 0.710 1.320 1.590 ;
        RECT  1.020 0.710 1.200 0.830 ;
        RECT  0.635 1.400 1.200 1.520 ;
        RECT  0.205 0.470 0.255 0.855 ;
        RECT  0.205 1.710 0.255 1.880 ;
        RECT  0.085 0.470 0.205 1.880 ;
    END
END EDFFHQX4AD
MACRO EDFFHQX8AD
    CLASS CORE ;
    FOREIGN EDFFHQX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.785 0.370 14.955 2.120 ;
        RECT  14.210 1.005 14.785 1.515 ;
        RECT  14.090 0.340 14.210 2.165 ;
        END
        AntennaDiffArea 0.86 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.100 1.125 3.220 1.900 ;
        RECT  2.055 1.125 3.100 1.360 ;
        RECT  0.420 1.780 3.100 1.900 ;
        RECT  0.160 1.780 0.420 1.960 ;
        END
        AntennaGateArea 0.269 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.055 1.325 1.225 ;
        RECT  0.580 0.910 0.830 1.225 ;
        END
        AntennaGateArea 0.49 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.225 0.910 4.655 1.170 ;
        END
        AntennaGateArea 0.281 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.315 -0.210 15.400 0.210 ;
        RECT  15.145 -0.210 15.315 0.800 ;
        RECT  14.595 -0.210 15.145 0.210 ;
        RECT  14.425 -0.210 14.595 0.800 ;
        RECT  13.865 -0.210 14.425 0.210 ;
        RECT  13.695 -0.210 13.865 0.525 ;
        RECT  12.660 -0.210 13.695 0.210 ;
        RECT  12.140 -0.210 12.660 0.255 ;
        RECT  9.945 -0.210 12.140 0.210 ;
        RECT  9.685 -0.210 9.945 0.260 ;
        RECT  9.165 -0.210 9.685 0.210 ;
        RECT  8.905 -0.210 9.165 0.260 ;
        RECT  7.820 -0.210 8.905 0.210 ;
        RECT  7.300 -0.210 7.820 0.260 ;
        RECT  5.755 -0.210 7.300 0.210 ;
        RECT  5.495 -0.210 5.755 0.260 ;
        RECT  4.560 -0.210 5.495 0.210 ;
        RECT  4.300 -0.210 4.560 0.255 ;
        RECT  3.860 -0.210 4.300 0.210 ;
        RECT  3.600 -0.210 3.860 0.300 ;
        RECT  1.785 -0.210 3.600 0.210 ;
        RECT  1.525 -0.210 1.785 0.260 ;
        RECT  0.920 -0.210 1.525 0.210 ;
        RECT  0.400 -0.210 0.920 0.330 ;
        RECT  0.000 -0.210 0.400 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.290 2.310 15.400 2.730 ;
        RECT  15.170 1.635 15.290 2.730 ;
        RECT  14.595 2.310 15.170 2.730 ;
        RECT  14.425 1.680 14.595 2.730 ;
        RECT  13.865 2.310 14.425 2.730 ;
        RECT  13.695 1.795 13.865 2.730 ;
        RECT  13.315 2.310 13.695 2.730 ;
        RECT  13.145 1.950 13.315 2.730 ;
        RECT  10.300 2.310 13.145 2.730 ;
        RECT  10.040 2.260 10.300 2.730 ;
        RECT  9.540 2.310 10.040 2.730 ;
        RECT  9.280 2.260 9.540 2.730 ;
        RECT  8.760 2.310 9.280 2.730 ;
        RECT  8.500 2.260 8.760 2.730 ;
        RECT  6.540 2.310 8.500 2.730 ;
        RECT  6.020 2.260 6.540 2.730 ;
        RECT  5.425 2.310 6.020 2.730 ;
        RECT  5.165 2.260 5.425 2.730 ;
        RECT  3.815 2.310 5.165 2.730 ;
        RECT  3.645 1.995 3.815 2.730 ;
        RECT  2.005 2.310 3.645 2.730 ;
        RECT  1.835 2.050 2.005 2.730 ;
        RECT  1.285 2.310 1.835 2.730 ;
        RECT  1.115 2.045 1.285 2.730 ;
        RECT  0.565 2.310 1.115 2.730 ;
        RECT  0.395 2.090 0.565 2.730 ;
        RECT  0.000 2.310 0.395 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 15.400 2.520 ;
        LAYER M1 ;
        RECT  13.845 0.735 13.965 1.600 ;
        RECT  13.410 0.735 13.845 0.880 ;
        RECT  13.435 1.430 13.845 1.600 ;
        RECT  12.860 1.005 13.725 1.265 ;
        RECT  13.315 1.430 13.435 1.780 ;
        RECT  13.265 0.380 13.410 0.880 ;
        RECT  12.930 1.660 13.315 1.780 ;
        RECT  4.390 0.380 13.265 0.500 ;
        RECT  12.810 1.660 12.930 2.090 ;
        RECT  12.740 0.620 12.860 1.540 ;
        RECT  10.425 0.620 12.740 0.740 ;
        RECT  12.435 1.420 12.740 1.540 ;
        RECT  7.775 2.020 12.670 2.140 ;
        RECT  12.475 1.140 12.615 1.260 ;
        RECT  12.355 0.950 12.475 1.260 ;
        RECT  12.430 1.420 12.435 1.850 ;
        RECT  12.260 1.420 12.430 1.900 ;
        RECT  11.335 0.950 12.355 1.070 ;
        RECT  10.780 1.780 12.260 1.900 ;
        RECT  11.070 1.540 12.120 1.660 ;
        RECT  10.950 0.860 11.070 1.660 ;
        RECT  10.255 0.860 10.950 0.980 ;
        RECT  10.635 1.530 10.950 1.660 ;
        RECT  10.015 1.120 10.805 1.240 ;
        RECT  10.465 1.530 10.635 1.800 ;
        RECT  9.775 1.680 10.465 1.800 ;
        RECT  10.135 0.720 10.255 0.980 ;
        RECT  9.895 0.620 10.015 1.240 ;
        RECT  8.695 0.620 9.895 0.740 ;
        RECT  9.655 0.860 9.775 1.800 ;
        RECT  9.285 0.860 9.655 0.980 ;
        RECT  8.520 1.680 9.655 1.800 ;
        RECT  9.030 1.185 9.460 1.355 ;
        RECT  8.910 1.000 9.030 1.355 ;
        RECT  8.280 1.000 8.910 1.120 ;
        RECT  8.435 0.620 8.695 0.780 ;
        RECT  8.400 1.305 8.520 1.800 ;
        RECT  5.810 0.620 8.435 0.740 ;
        RECT  8.160 1.000 8.280 1.550 ;
        RECT  8.065 1.430 8.160 1.550 ;
        RECT  7.895 1.430 8.065 1.840 ;
        RECT  7.275 1.430 7.895 1.550 ;
        RECT  7.655 1.685 7.775 2.140 ;
        RECT  6.810 0.965 7.670 1.085 ;
        RECT  6.810 1.685 7.655 1.805 ;
        RECT  7.355 1.930 7.475 2.190 ;
        RECT  4.115 2.020 7.355 2.140 ;
        RECT  7.105 1.320 7.275 1.550 ;
        RECT  6.690 0.965 6.810 1.805 ;
        RECT  5.815 1.685 6.690 1.805 ;
        RECT  5.695 1.685 5.815 1.900 ;
        RECT  5.690 0.620 5.810 1.520 ;
        RECT  4.470 1.780 5.695 1.900 ;
        RECT  5.110 0.620 5.690 0.780 ;
        RECT  5.375 1.400 5.690 1.520 ;
        RECT  5.135 0.965 5.570 1.135 ;
        RECT  5.255 1.400 5.375 1.660 ;
        RECT  4.755 1.540 5.255 1.660 ;
        RECT  4.990 0.965 5.135 1.420 ;
        RECT  4.875 0.640 4.990 1.420 ;
        RECT  4.825 0.640 4.875 1.135 ;
        RECT  4.730 0.640 4.825 0.760 ;
        RECT  4.635 1.400 4.755 1.660 ;
        RECT  4.350 1.495 4.470 1.900 ;
        RECT  4.270 0.380 4.390 0.540 ;
        RECT  4.080 1.495 4.350 1.615 ;
        RECT  3.700 0.420 4.270 0.540 ;
        RECT  4.080 0.660 4.240 0.780 ;
        RECT  3.995 1.735 4.115 2.140 ;
        RECT  3.960 0.660 4.080 1.615 ;
        RECT  3.460 1.735 3.995 1.855 ;
        RECT  3.580 0.420 3.700 1.190 ;
        RECT  3.340 0.620 3.460 2.140 ;
        RECT  1.815 0.620 3.340 0.740 ;
        RECT  2.130 2.020 3.340 2.140 ;
        RECT  2.775 0.330 3.035 0.500 ;
        RECT  1.585 0.380 2.775 0.500 ;
        RECT  1.695 1.540 2.750 1.660 ;
        RECT  1.695 0.860 2.455 0.980 ;
        RECT  1.575 0.710 1.695 1.660 ;
        RECT  1.465 0.380 1.585 0.590 ;
        RECT  1.095 0.710 1.575 0.830 ;
        RECT  0.710 1.540 1.575 1.660 ;
        RECT  0.230 0.470 1.465 0.590 ;
        RECT  0.110 0.470 0.230 1.625 ;
    END
END EDFFHQX8AD
MACRO EDFFTRX1AD
    CLASS CORE ;
    FOREIGN EDFFTRX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.910 1.870 1.070 ;
        END
        AntennaGateArea 0.04 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.470 0.685 8.610 1.910 ;
        RECT  8.425 0.685 8.470 0.855 ;
        RECT  8.440 1.390 8.470 1.910 ;
        END
        AntennaDiffArea 0.207 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.860 1.145 8.065 1.375 ;
        RECT  7.855 0.640 7.860 1.375 ;
        RECT  7.690 0.640 7.855 1.610 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.110 2.540 1.310 ;
        RECT  1.210 1.190 2.280 1.310 ;
        RECT  1.090 1.190 1.210 1.685 ;
        RECT  0.490 1.565 1.090 1.685 ;
        RECT  0.350 0.980 0.490 1.685 ;
        END
        AntennaGateArea 0.088 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.990 1.965 2.170 ;
        END
        AntennaGateArea 0.04 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.900 1.230 1.070 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.235 -0.210 8.680 0.210 ;
        RECT  8.065 -0.210 8.235 0.855 ;
        RECT  7.150 -0.210 8.065 0.210 ;
        RECT  6.890 -0.210 7.150 0.520 ;
        RECT  5.825 -0.210 6.890 0.210 ;
        RECT  5.705 -0.210 5.825 0.800 ;
        RECT  4.500 -0.210 5.705 0.210 ;
        RECT  4.240 -0.210 4.500 0.695 ;
        RECT  1.305 -0.210 4.240 0.210 ;
        RECT  1.135 -0.210 1.305 0.540 ;
        RECT  0.585 -0.210 1.135 0.210 ;
        RECT  0.415 -0.210 0.585 0.395 ;
        RECT  0.000 -0.210 0.415 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.215 2.310 8.680 2.730 ;
        RECT  8.045 1.970 8.215 2.730 ;
        RECT  7.150 2.310 8.045 2.730 ;
        RECT  7.010 1.910 7.150 2.730 ;
        RECT  5.610 2.310 7.010 2.730 ;
        RECT  5.350 2.240 5.610 2.730 ;
        RECT  4.505 2.310 5.350 2.730 ;
        RECT  4.245 2.240 4.505 2.730 ;
        RECT  2.415 2.310 4.245 2.730 ;
        RECT  2.245 2.125 2.415 2.730 ;
        RECT  1.305 2.310 2.245 2.730 ;
        RECT  1.135 2.045 1.305 2.730 ;
        RECT  0.575 2.310 1.135 2.730 ;
        RECT  0.405 2.045 0.575 2.730 ;
        RECT  0.000 2.310 0.405 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.680 2.520 ;
        LAYER M1 ;
        RECT  8.305 1.010 8.330 1.270 ;
        RECT  8.185 1.010 8.305 1.850 ;
        RECT  7.565 1.730 8.185 1.850 ;
        RECT  7.445 0.685 7.565 1.850 ;
        RECT  7.325 0.685 7.445 0.855 ;
        RECT  6.890 1.485 7.445 1.655 ;
        RECT  7.200 1.005 7.320 1.265 ;
        RECT  7.005 1.005 7.200 1.125 ;
        RECT  6.885 0.640 7.005 1.125 ;
        RECT  6.750 1.485 6.890 2.120 ;
        RECT  6.305 0.640 6.885 0.760 ;
        RECT  6.630 1.980 6.750 2.120 ;
        RECT  6.510 0.880 6.630 1.860 ;
        RECT  2.655 2.000 6.630 2.120 ;
        RECT  6.450 0.880 6.510 1.140 ;
        RECT  3.525 1.740 6.510 1.860 ;
        RECT  6.065 0.330 6.400 0.450 ;
        RECT  6.305 1.445 6.355 1.615 ;
        RECT  6.185 0.640 6.305 1.615 ;
        RECT  5.945 0.330 6.065 1.595 ;
        RECT  5.335 1.425 5.945 1.595 ;
        RECT  5.680 0.920 5.800 1.180 ;
        RECT  5.585 0.920 5.680 1.040 ;
        RECT  5.465 0.405 5.585 1.040 ;
        RECT  4.890 0.405 5.465 0.525 ;
        RECT  5.165 0.665 5.335 1.595 ;
        RECT  5.015 1.425 5.165 1.595 ;
        RECT  4.770 0.405 4.890 1.490 ;
        RECT  4.710 0.405 4.770 0.810 ;
        RECT  4.350 1.370 4.770 1.490 ;
        RECT  4.590 0.930 4.620 1.190 ;
        RECT  4.470 0.815 4.590 1.190 ;
        RECT  3.815 0.815 4.470 0.935 ;
        RECT  4.230 1.055 4.350 1.490 ;
        RECT  4.090 1.055 4.230 1.175 ;
        RECT  3.645 0.620 3.815 1.505 ;
        RECT  3.485 0.620 3.645 0.740 ;
        RECT  3.405 0.965 3.525 1.860 ;
        RECT  3.270 0.965 3.405 1.085 ;
        RECT  3.165 1.290 3.285 1.865 ;
        RECT  3.150 0.860 3.270 1.085 ;
        RECT  1.775 1.720 3.165 1.865 ;
        RECT  2.270 0.860 3.150 0.980 ;
        RECT  2.680 1.100 2.800 1.560 ;
        RECT  1.450 1.440 2.680 1.560 ;
        RECT  2.520 0.620 2.660 0.740 ;
        RECT  2.400 0.420 2.520 0.740 ;
        RECT  1.490 0.420 2.400 0.540 ;
        RECT  2.150 0.660 2.270 0.980 ;
        RECT  0.925 0.660 2.150 0.780 ;
        RECT  1.605 1.695 1.775 1.865 ;
        RECT  1.330 1.440 1.450 1.925 ;
        RECT  0.230 1.805 1.330 1.925 ;
        RECT  0.740 1.325 0.970 1.445 ;
        RECT  0.755 0.540 0.925 0.780 ;
        RECT  0.740 0.660 0.755 0.780 ;
        RECT  0.620 0.660 0.740 1.445 ;
        RECT  0.090 0.610 0.230 1.925 ;
    END
END EDFFTRX1AD
MACRO EDFFTRX2AD
    CLASS CORE ;
    FOREIGN EDFFTRX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.910 1.870 1.070 ;
        END
        AntennaGateArea 0.04 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.470 0.330 8.610 2.190 ;
        RECT  8.440 0.330 8.470 0.850 ;
        RECT  8.440 1.410 8.470 2.190 ;
        END
        AntennaDiffArea 0.373 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.875 1.145 8.050 1.375 ;
        RECT  7.860 1.145 7.875 1.610 ;
        RECT  7.690 0.330 7.860 1.610 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.110 2.540 1.310 ;
        RECT  1.210 1.190 2.280 1.310 ;
        RECT  1.090 1.190 1.210 1.685 ;
        RECT  0.490 1.565 1.090 1.685 ;
        RECT  0.350 0.980 0.490 1.685 ;
        END
        AntennaGateArea 0.088 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.580 2.015 1.965 2.185 ;
        END
        AntennaGateArea 0.04 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.900 1.230 1.070 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.235 -0.210 8.680 0.210 ;
        RECT  8.065 -0.210 8.235 0.805 ;
        RECT  7.200 -0.210 8.065 0.210 ;
        RECT  6.940 -0.210 7.200 0.520 ;
        RECT  5.825 -0.210 6.940 0.210 ;
        RECT  5.705 -0.210 5.825 0.800 ;
        RECT  4.500 -0.210 5.705 0.210 ;
        RECT  4.240 -0.210 4.500 0.695 ;
        RECT  1.305 -0.210 4.240 0.210 ;
        RECT  1.135 -0.210 1.305 0.540 ;
        RECT  0.585 -0.210 1.135 0.210 ;
        RECT  0.415 -0.210 0.585 0.395 ;
        RECT  0.000 -0.210 0.415 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.235 2.310 8.680 2.730 ;
        RECT  8.065 1.970 8.235 2.730 ;
        RECT  7.205 2.310 8.065 2.730 ;
        RECT  7.065 2.010 7.205 2.730 ;
        RECT  5.610 2.310 7.065 2.730 ;
        RECT  5.350 2.240 5.610 2.730 ;
        RECT  4.505 2.310 5.350 2.730 ;
        RECT  4.245 2.240 4.505 2.730 ;
        RECT  2.415 2.310 4.245 2.730 ;
        RECT  2.245 2.145 2.415 2.730 ;
        RECT  1.305 2.310 2.245 2.730 ;
        RECT  1.135 2.045 1.305 2.730 ;
        RECT  0.575 2.310 1.135 2.730 ;
        RECT  0.405 2.045 0.575 2.730 ;
        RECT  0.000 2.310 0.405 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.680 2.520 ;
        LAYER M1 ;
        RECT  8.305 1.010 8.350 1.270 ;
        RECT  8.185 1.010 8.305 1.850 ;
        RECT  7.565 1.730 8.185 1.850 ;
        RECT  7.445 0.680 7.565 1.850 ;
        RECT  7.365 0.680 7.445 0.850 ;
        RECT  6.945 1.550 7.445 1.720 ;
        RECT  7.200 1.005 7.320 1.265 ;
        RECT  7.005 1.005 7.200 1.125 ;
        RECT  6.885 0.640 7.005 1.125 ;
        RECT  6.805 1.550 6.945 2.140 ;
        RECT  6.305 0.640 6.885 0.760 ;
        RECT  5.850 2.020 6.805 2.140 ;
        RECT  6.565 0.930 6.685 1.900 ;
        RECT  6.500 0.930 6.565 1.190 ;
        RECT  6.090 1.780 6.565 1.900 ;
        RECT  6.305 1.520 6.445 1.640 ;
        RECT  6.065 0.330 6.400 0.450 ;
        RECT  6.185 0.640 6.305 1.640 ;
        RECT  5.970 1.760 6.090 1.900 ;
        RECT  5.945 0.330 6.065 1.595 ;
        RECT  3.525 1.760 5.970 1.880 ;
        RECT  5.335 1.425 5.945 1.595 ;
        RECT  5.730 2.000 5.850 2.140 ;
        RECT  5.680 0.920 5.800 1.250 ;
        RECT  2.915 2.000 5.730 2.120 ;
        RECT  5.585 0.920 5.680 1.040 ;
        RECT  5.465 0.405 5.585 1.040 ;
        RECT  4.890 0.405 5.465 0.525 ;
        RECT  5.185 0.665 5.335 1.595 ;
        RECT  5.165 0.665 5.185 1.620 ;
        RECT  5.015 1.425 5.165 1.620 ;
        RECT  4.770 0.405 4.890 1.490 ;
        RECT  4.710 0.405 4.770 0.810 ;
        RECT  4.350 1.370 4.770 1.490 ;
        RECT  4.590 0.930 4.620 1.190 ;
        RECT  4.470 0.815 4.590 1.190 ;
        RECT  3.815 0.815 4.470 0.935 ;
        RECT  4.230 1.055 4.350 1.490 ;
        RECT  4.090 1.055 4.230 1.175 ;
        RECT  3.645 0.620 3.815 1.505 ;
        RECT  3.485 0.620 3.645 0.740 ;
        RECT  3.405 0.965 3.525 1.880 ;
        RECT  3.270 0.965 3.405 1.085 ;
        RECT  3.165 1.290 3.285 1.865 ;
        RECT  3.150 0.860 3.270 1.085 ;
        RECT  1.775 1.715 3.165 1.865 ;
        RECT  2.270 0.860 3.150 0.980 ;
        RECT  2.655 2.000 2.915 2.150 ;
        RECT  2.680 1.100 2.800 1.550 ;
        RECT  1.450 1.430 2.680 1.550 ;
        RECT  2.520 0.620 2.660 0.740 ;
        RECT  2.400 0.420 2.520 0.740 ;
        RECT  1.490 0.420 2.400 0.540 ;
        RECT  2.150 0.660 2.270 0.980 ;
        RECT  0.925 0.660 2.150 0.780 ;
        RECT  1.605 1.715 1.775 1.895 ;
        RECT  1.330 1.430 1.450 1.925 ;
        RECT  0.230 1.805 1.330 1.925 ;
        RECT  0.740 1.325 0.970 1.445 ;
        RECT  0.755 0.540 0.925 0.780 ;
        RECT  0.740 0.660 0.755 0.780 ;
        RECT  0.620 0.660 0.740 1.445 ;
        RECT  0.090 0.610 0.230 1.925 ;
    END
END EDFFTRX2AD
MACRO EDFFTRX4AD
    CLASS CORE ;
    FOREIGN EDFFTRX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.910 1.870 1.070 ;
        END
        AntennaGateArea 0.04 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.635 0.365 9.730 1.795 ;
        RECT  9.590 0.365 9.635 2.170 ;
        RECT  9.465 0.365 9.590 0.795 ;
        RECT  9.465 1.480 9.590 2.170 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.720 0.410 8.890 1.640 ;
        END
        AntennaDiffArea 0.454 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.325 1.110 2.495 1.310 ;
        RECT  1.200 1.190 2.325 1.310 ;
        RECT  1.080 1.190 1.200 1.685 ;
        RECT  0.490 1.565 1.080 1.685 ;
        RECT  0.350 0.975 0.490 1.685 ;
        END
        AntennaGateArea 0.088 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 2.005 1.965 2.170 ;
        END
        AntennaGateArea 0.04 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.900 1.230 1.070 ;
        END
        AntennaGateArea 0.096 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.970 -0.210 10.080 0.210 ;
        RECT  9.850 -0.210 9.970 0.840 ;
        RECT  9.270 -0.210 9.850 0.210 ;
        RECT  9.100 -0.210 9.270 0.795 ;
        RECT  8.520 -0.210 9.100 0.210 ;
        RECT  8.350 -0.210 8.520 0.675 ;
        RECT  7.820 -0.210 8.350 0.210 ;
        RECT  7.650 -0.210 7.820 0.810 ;
        RECT  6.920 -0.210 7.650 0.210 ;
        RECT  6.660 -0.210 6.920 0.300 ;
        RECT  5.660 -0.210 6.660 0.210 ;
        RECT  5.400 -0.210 5.660 0.300 ;
        RECT  4.490 -0.210 5.400 0.210 ;
        RECT  4.230 -0.210 4.490 0.650 ;
        RECT  1.350 -0.210 4.230 0.210 ;
        RECT  1.090 -0.210 1.350 0.540 ;
        RECT  0.585 -0.210 1.090 0.210 ;
        RECT  0.415 -0.210 0.585 0.395 ;
        RECT  0.000 -0.210 0.415 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.970 2.310 10.080 2.730 ;
        RECT  9.850 1.435 9.970 2.730 ;
        RECT  9.260 2.310 9.850 2.730 ;
        RECT  9.090 2.010 9.260 2.730 ;
        RECT  8.520 2.310 9.090 2.730 ;
        RECT  8.350 2.010 8.520 2.730 ;
        RECT  7.845 2.310 8.350 2.730 ;
        RECT  7.585 2.220 7.845 2.730 ;
        RECT  6.920 2.310 7.585 2.730 ;
        RECT  6.660 2.220 6.920 2.730 ;
        RECT  5.655 2.310 6.660 2.730 ;
        RECT  5.395 2.220 5.655 2.730 ;
        RECT  4.500 2.310 5.395 2.730 ;
        RECT  4.240 2.220 4.500 2.730 ;
        RECT  2.390 2.310 4.240 2.730 ;
        RECT  2.220 2.135 2.390 2.730 ;
        RECT  1.315 2.310 2.220 2.730 ;
        RECT  1.145 2.045 1.315 2.730 ;
        RECT  0.575 2.310 1.145 2.730 ;
        RECT  0.405 2.045 0.575 2.730 ;
        RECT  0.000 2.310 0.405 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.080 2.520 ;
        LAYER M1 ;
        RECT  9.290 1.010 9.460 1.270 ;
        RECT  9.170 1.010 9.290 1.890 ;
        RECT  8.590 1.770 9.170 1.890 ;
        RECT  8.470 0.795 8.590 1.890 ;
        RECT  8.180 0.795 8.470 0.915 ;
        RECT  8.155 1.770 8.470 1.890 ;
        RECT  7.520 1.055 8.320 1.225 ;
        RECT  8.010 0.640 8.180 0.915 ;
        RECT  8.035 1.370 8.155 2.100 ;
        RECT  2.870 1.980 8.035 2.100 ;
        RECT  7.400 0.610 7.520 1.615 ;
        RECT  7.170 0.610 7.400 0.730 ;
        RECT  7.060 1.495 7.400 1.615 ;
        RECT  7.160 0.850 7.280 1.360 ;
        RECT  7.000 0.545 7.170 0.730 ;
        RECT  6.180 0.850 7.160 0.970 ;
        RECT  6.940 1.495 7.060 1.860 ;
        RECT  6.030 0.610 7.000 0.730 ;
        RECT  6.805 1.090 6.975 1.365 ;
        RECT  6.030 1.740 6.940 1.860 ;
        RECT  6.370 1.245 6.805 1.365 ;
        RECT  6.250 1.245 6.370 1.615 ;
        RECT  5.765 1.495 6.250 1.615 ;
        RECT  6.040 0.850 6.180 1.125 ;
        RECT  5.920 0.850 6.040 1.375 ;
        RECT  5.230 1.255 5.920 1.375 ;
        RECT  5.695 0.995 5.800 1.135 ;
        RECT  5.645 1.495 5.765 1.860 ;
        RECT  5.540 0.420 5.695 1.135 ;
        RECT  3.525 1.740 5.645 1.860 ;
        RECT  4.875 0.420 5.540 0.540 ;
        RECT  5.115 0.660 5.320 0.780 ;
        RECT  5.115 1.255 5.230 1.595 ;
        RECT  4.995 0.660 5.115 1.595 ;
        RECT  4.755 0.420 4.875 1.515 ;
        RECT  4.695 0.420 4.755 0.795 ;
        RECT  4.675 1.345 4.755 1.515 ;
        RECT  4.280 1.345 4.675 1.465 ;
        RECT  4.575 0.915 4.635 1.175 ;
        RECT  4.455 0.770 4.575 1.175 ;
        RECT  3.790 0.770 4.455 0.890 ;
        RECT  4.160 1.010 4.280 1.465 ;
        RECT  3.670 0.630 3.790 1.550 ;
        RECT  3.485 0.630 3.670 0.750 ;
        RECT  3.405 0.870 3.525 1.860 ;
        RECT  3.150 0.870 3.405 1.085 ;
        RECT  3.165 1.290 3.285 1.850 ;
        RECT  1.730 1.705 3.165 1.850 ;
        RECT  2.270 0.870 3.150 0.990 ;
        RECT  2.700 1.980 2.870 2.185 ;
        RECT  2.655 1.110 2.825 1.570 ;
        RECT  2.520 0.630 2.660 0.750 ;
        RECT  1.440 1.450 2.655 1.570 ;
        RECT  2.400 0.420 2.520 0.750 ;
        RECT  1.490 0.420 2.400 0.540 ;
        RECT  2.150 0.660 2.270 0.990 ;
        RECT  0.925 0.660 2.150 0.780 ;
        RECT  1.560 1.705 1.730 1.875 ;
        RECT  1.320 1.450 1.440 1.925 ;
        RECT  0.230 1.805 1.320 1.925 ;
        RECT  0.740 1.325 0.960 1.445 ;
        RECT  0.740 0.540 0.925 0.780 ;
        RECT  0.620 0.540 0.740 1.445 ;
        RECT  0.090 0.610 0.230 1.925 ;
    END
END EDFFTRX4AD
MACRO EDFFTRXLAD
    CLASS CORE ;
    FOREIGN EDFFTRXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.910 1.870 1.070 ;
        END
        AntennaGateArea 0.04 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.470 0.720 8.610 1.640 ;
        RECT  8.425 0.720 8.470 0.890 ;
        RECT  8.425 1.470 8.470 1.640 ;
        END
        AntennaDiffArea 0.143 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.860 1.145 8.065 1.375 ;
        RECT  7.855 0.675 7.860 1.375 ;
        RECT  7.690 0.675 7.855 1.610 ;
        END
        AntennaDiffArea 0.143 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.110 2.540 1.310 ;
        RECT  1.210 1.190 2.280 1.310 ;
        RECT  1.090 1.190 1.210 1.685 ;
        RECT  0.490 1.565 1.090 1.685 ;
        RECT  0.350 0.980 0.490 1.685 ;
        END
        AntennaGateArea 0.088 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.990 1.965 2.170 ;
        END
        AntennaGateArea 0.04 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.900 1.230 1.070 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.235 -0.210 8.680 0.210 ;
        RECT  8.065 -0.210 8.235 0.890 ;
        RECT  7.150 -0.210 8.065 0.210 ;
        RECT  6.890 -0.210 7.150 0.520 ;
        RECT  5.815 -0.210 6.890 0.210 ;
        RECT  5.695 -0.210 5.815 0.800 ;
        RECT  4.500 -0.210 5.695 0.210 ;
        RECT  4.240 -0.210 4.500 0.695 ;
        RECT  1.305 -0.210 4.240 0.210 ;
        RECT  1.135 -0.210 1.305 0.540 ;
        RECT  0.585 -0.210 1.135 0.210 ;
        RECT  0.415 -0.210 0.585 0.395 ;
        RECT  0.000 -0.210 0.415 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.215 2.310 8.680 2.730 ;
        RECT  8.045 1.970 8.215 2.730 ;
        RECT  7.150 2.310 8.045 2.730 ;
        RECT  7.010 1.910 7.150 2.730 ;
        RECT  5.610 2.310 7.010 2.730 ;
        RECT  5.350 2.240 5.610 2.730 ;
        RECT  4.505 2.310 5.350 2.730 ;
        RECT  4.245 2.240 4.505 2.730 ;
        RECT  2.415 2.310 4.245 2.730 ;
        RECT  2.245 2.125 2.415 2.730 ;
        RECT  1.305 2.310 2.245 2.730 ;
        RECT  1.135 2.045 1.305 2.730 ;
        RECT  0.575 2.310 1.135 2.730 ;
        RECT  0.405 2.045 0.575 2.730 ;
        RECT  0.000 2.310 0.405 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.680 2.520 ;
        LAYER M1 ;
        RECT  8.305 1.010 8.330 1.270 ;
        RECT  8.185 1.010 8.305 1.850 ;
        RECT  7.565 1.730 8.185 1.850 ;
        RECT  7.445 0.685 7.565 1.850 ;
        RECT  7.325 0.685 7.445 0.855 ;
        RECT  6.890 1.485 7.445 1.655 ;
        RECT  7.200 1.005 7.320 1.265 ;
        RECT  7.005 1.005 7.200 1.125 ;
        RECT  6.885 0.640 7.005 1.125 ;
        RECT  6.750 1.485 6.890 2.120 ;
        RECT  6.305 0.640 6.885 0.760 ;
        RECT  2.655 2.000 6.750 2.120 ;
        RECT  6.510 0.880 6.630 1.860 ;
        RECT  6.450 0.880 6.510 1.140 ;
        RECT  3.525 1.740 6.510 1.860 ;
        RECT  6.065 0.330 6.400 0.450 ;
        RECT  6.305 1.445 6.355 1.615 ;
        RECT  6.185 0.640 6.305 1.615 ;
        RECT  5.945 0.330 6.065 1.595 ;
        RECT  5.335 1.425 5.945 1.595 ;
        RECT  5.680 0.920 5.800 1.180 ;
        RECT  5.575 0.920 5.680 1.040 ;
        RECT  5.455 0.395 5.575 1.040 ;
        RECT  4.890 0.395 5.455 0.515 ;
        RECT  5.165 0.635 5.335 1.595 ;
        RECT  5.015 1.425 5.165 1.595 ;
        RECT  4.770 0.395 4.890 1.490 ;
        RECT  4.710 0.395 4.770 0.810 ;
        RECT  4.350 1.370 4.770 1.490 ;
        RECT  4.590 0.930 4.620 1.190 ;
        RECT  4.470 0.815 4.590 1.190 ;
        RECT  3.815 0.815 4.470 0.935 ;
        RECT  4.230 1.055 4.350 1.490 ;
        RECT  4.090 1.055 4.230 1.175 ;
        RECT  3.645 0.620 3.815 1.505 ;
        RECT  3.485 0.620 3.645 0.740 ;
        RECT  3.405 0.965 3.525 1.860 ;
        RECT  3.270 0.965 3.405 1.085 ;
        RECT  3.165 1.290 3.285 1.865 ;
        RECT  3.150 0.860 3.270 1.085 ;
        RECT  1.775 1.720 3.165 1.865 ;
        RECT  2.270 0.860 3.150 0.980 ;
        RECT  2.680 1.100 2.800 1.560 ;
        RECT  1.450 1.440 2.680 1.560 ;
        RECT  2.520 0.620 2.660 0.740 ;
        RECT  2.400 0.420 2.520 0.740 ;
        RECT  1.490 0.420 2.400 0.540 ;
        RECT  2.150 0.660 2.270 0.980 ;
        RECT  0.925 0.660 2.150 0.780 ;
        RECT  1.605 1.695 1.775 1.865 ;
        RECT  1.330 1.440 1.450 1.925 ;
        RECT  0.230 1.805 1.330 1.925 ;
        RECT  0.740 1.325 0.970 1.445 ;
        RECT  0.755 0.540 0.925 0.780 ;
        RECT  0.740 0.660 0.755 0.780 ;
        RECT  0.620 0.660 0.740 1.445 ;
        RECT  0.090 0.610 0.230 1.925 ;
    END
END EDFFTRXLAD
MACRO EDFFX1AD
    CLASS CORE ;
    FOREIGN EDFFX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 1.425 7.490 1.920 ;
        RECT  7.330 0.625 7.450 1.920 ;
        END
        AntennaDiffArea 0.207 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.865 6.970 1.860 ;
        RECT  6.730 0.865 6.850 1.095 ;
        RECT  6.260 1.740 6.850 1.860 ;
        RECT  6.610 0.605 6.730 1.095 ;
        END
        AntennaDiffArea 0.183 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.170 0.910 0.570 1.095 ;
        END
        AntennaGateArea 0.119 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.930 0.865 1.375 1.050 ;
        END
        AntennaGateArea 0.071 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.100 1.130 3.455 1.355 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.160 -0.210 7.560 0.210 ;
        RECT  6.900 -0.210 7.160 0.745 ;
        RECT  6.140 -0.210 6.900 0.210 ;
        RECT  5.880 -0.210 6.140 0.445 ;
        RECT  4.685 -0.210 5.880 0.210 ;
        RECT  4.425 -0.210 4.685 0.415 ;
        RECT  3.470 -0.210 4.425 0.210 ;
        RECT  3.210 -0.210 3.470 0.415 ;
        RECT  1.575 -0.210 3.210 0.210 ;
        RECT  1.405 -0.210 1.575 0.260 ;
        RECT  0.545 -0.210 1.405 0.210 ;
        RECT  0.375 -0.210 0.545 0.335 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.140 2.310 7.560 2.730 ;
        RECT  6.880 2.220 7.140 2.730 ;
        RECT  6.140 2.310 6.880 2.730 ;
        RECT  5.880 2.220 6.140 2.730 ;
        RECT  4.890 2.310 5.880 2.730 ;
        RECT  4.630 2.220 4.890 2.730 ;
        RECT  3.780 2.310 4.630 2.730 ;
        RECT  3.520 2.220 3.780 2.730 ;
        RECT  3.060 2.310 3.520 2.730 ;
        RECT  2.800 2.250 3.060 2.730 ;
        RECT  1.425 2.310 2.800 2.730 ;
        RECT  1.255 1.720 1.425 2.730 ;
        RECT  0.610 2.310 1.255 2.730 ;
        RECT  0.490 2.055 0.610 2.730 ;
        RECT  0.000 2.310 0.490 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  7.090 1.005 7.210 2.100 ;
        RECT  5.900 1.980 7.090 2.100 ;
        RECT  6.610 1.330 6.730 1.590 ;
        RECT  6.490 1.330 6.610 1.450 ;
        RECT  6.370 0.755 6.490 1.450 ;
        RECT  6.170 0.755 6.370 0.875 ;
        RECT  5.900 1.330 6.370 1.450 ;
        RECT  6.080 1.000 6.250 1.210 ;
        RECT  5.640 1.000 6.080 1.120 ;
        RECT  5.780 1.300 5.900 2.100 ;
        RECT  2.590 1.980 5.780 2.100 ;
        RECT  5.520 0.755 5.640 1.800 ;
        RECT  5.360 0.375 5.620 0.570 ;
        RECT  5.290 0.755 5.520 1.015 ;
        RECT  5.260 1.680 5.520 1.800 ;
        RECT  5.170 1.385 5.400 1.520 ;
        RECT  5.170 0.450 5.360 0.570 ;
        RECT  5.050 0.450 5.170 1.520 ;
        RECT  4.750 1.085 5.050 1.205 ;
        RECT  4.805 0.375 4.925 0.655 ;
        RECT  4.020 0.535 4.805 0.655 ;
        RECT  4.630 1.085 4.750 1.860 ;
        RECT  4.510 1.085 4.630 1.345 ;
        RECT  2.720 1.740 4.630 1.860 ;
        RECT  4.380 1.500 4.510 1.620 ;
        RECT  4.250 0.810 4.380 1.620 ;
        RECT  4.210 0.810 4.250 1.320 ;
        RECT  4.140 1.060 4.210 1.320 ;
        RECT  4.020 1.500 4.130 1.620 ;
        RECT  3.900 0.535 4.020 1.620 ;
        RECT  3.815 0.535 3.900 0.995 ;
        RECT  2.980 1.500 3.900 1.620 ;
        RECT  3.695 1.120 3.780 1.380 ;
        RECT  3.575 0.620 3.695 1.380 ;
        RECT  2.580 0.620 3.575 0.740 ;
        RECT  3.030 0.860 3.290 1.005 ;
        RECT  2.720 0.860 3.030 0.980 ;
        RECT  2.860 1.360 2.980 1.620 ;
        RECT  2.600 0.860 2.720 1.860 ;
        RECT  2.270 0.860 2.600 0.980 ;
        RECT  2.480 1.360 2.600 1.620 ;
        RECT  2.470 1.980 2.590 2.140 ;
        RECT  2.460 0.475 2.580 0.740 ;
        RECT  1.960 2.020 2.470 2.140 ;
        RECT  2.150 0.620 2.460 0.740 ;
        RECT  2.320 1.715 2.395 1.885 ;
        RECT  2.200 1.165 2.320 1.885 ;
        RECT  1.380 0.380 2.270 0.500 ;
        RECT  2.150 1.165 2.200 1.285 ;
        RECT  2.030 0.620 2.150 1.285 ;
        RECT  0.600 1.480 2.080 1.600 ;
        RECT  1.700 2.020 1.960 2.190 ;
        RECT  1.620 0.745 1.760 0.865 ;
        RECT  1.500 0.745 1.620 1.335 ;
        RECT  1.090 1.170 1.500 1.335 ;
        RECT  1.260 0.380 1.380 0.740 ;
        RECT  0.960 0.620 1.260 0.740 ;
        RECT  0.810 1.215 1.090 1.335 ;
        RECT  0.690 0.670 0.810 1.335 ;
        RECT  0.255 0.670 0.690 0.790 ;
        RECT  0.230 1.215 0.690 1.335 ;
        RECT  0.085 0.595 0.255 0.790 ;
        RECT  0.110 1.215 0.230 2.040 ;
    END
END EDFFX1AD
MACRO EDFFX2AD
    CLASS CORE ;
    FOREIGN EDFFX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 1.425 7.490 2.190 ;
        RECT  7.330 0.330 7.450 2.190 ;
        END
        AntennaDiffArea 0.373 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.865 6.970 1.860 ;
        RECT  6.730 0.865 6.850 1.095 ;
        RECT  6.260 1.740 6.850 1.860 ;
        RECT  6.610 0.330 6.730 1.095 ;
        END
        AntennaDiffArea 0.344 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.170 0.910 0.570 1.095 ;
        END
        AntennaGateArea 0.119 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.930 0.865 1.375 1.050 ;
        END
        AntennaGateArea 0.071 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.100 1.130 3.455 1.355 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.115 -0.210 7.560 0.210 ;
        RECT  6.945 -0.210 7.115 0.745 ;
        RECT  6.095 -0.210 6.945 0.210 ;
        RECT  5.925 -0.210 6.095 0.410 ;
        RECT  4.640 -0.210 5.925 0.210 ;
        RECT  4.380 -0.210 4.640 0.415 ;
        RECT  3.470 -0.210 4.380 0.210 ;
        RECT  3.210 -0.210 3.470 0.415 ;
        RECT  1.575 -0.210 3.210 0.210 ;
        RECT  1.405 -0.210 1.575 0.260 ;
        RECT  0.545 -0.210 1.405 0.210 ;
        RECT  0.375 -0.210 0.545 0.335 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.090 2.310 7.560 2.730 ;
        RECT  6.830 2.220 7.090 2.730 ;
        RECT  6.140 2.310 6.830 2.730 ;
        RECT  5.880 2.220 6.140 2.730 ;
        RECT  4.890 2.310 5.880 2.730 ;
        RECT  4.630 2.220 4.890 2.730 ;
        RECT  3.780 2.310 4.630 2.730 ;
        RECT  3.520 2.220 3.780 2.730 ;
        RECT  3.060 2.310 3.520 2.730 ;
        RECT  2.800 2.250 3.060 2.730 ;
        RECT  1.425 2.310 2.800 2.730 ;
        RECT  1.255 1.720 1.425 2.730 ;
        RECT  0.610 2.310 1.255 2.730 ;
        RECT  0.490 2.055 0.610 2.730 ;
        RECT  0.000 2.310 0.490 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  7.090 1.005 7.210 2.100 ;
        RECT  5.900 1.980 7.090 2.100 ;
        RECT  6.490 1.330 6.730 1.590 ;
        RECT  6.370 0.725 6.490 1.590 ;
        RECT  6.170 0.725 6.370 0.845 ;
        RECT  5.900 1.470 6.370 1.590 ;
        RECT  6.130 1.000 6.250 1.260 ;
        RECT  5.640 1.000 6.130 1.120 ;
        RECT  5.780 1.300 5.900 2.100 ;
        RECT  2.590 1.980 5.780 2.100 ;
        RECT  5.520 0.755 5.640 1.800 ;
        RECT  5.360 0.375 5.620 0.570 ;
        RECT  5.290 0.755 5.520 1.015 ;
        RECT  5.260 1.680 5.520 1.800 ;
        RECT  5.170 1.385 5.400 1.520 ;
        RECT  5.170 0.450 5.360 0.570 ;
        RECT  5.050 0.450 5.170 1.520 ;
        RECT  4.750 1.120 5.050 1.240 ;
        RECT  4.760 0.335 4.930 0.655 ;
        RECT  4.020 0.535 4.760 0.655 ;
        RECT  4.630 1.120 4.750 1.860 ;
        RECT  4.510 1.120 4.630 1.380 ;
        RECT  2.720 1.740 4.630 1.860 ;
        RECT  4.380 1.500 4.510 1.620 ;
        RECT  4.250 0.835 4.380 1.620 ;
        RECT  4.210 0.835 4.250 1.320 ;
        RECT  4.140 1.060 4.210 1.320 ;
        RECT  4.020 1.500 4.130 1.620 ;
        RECT  3.900 0.535 4.020 1.620 ;
        RECT  3.815 0.535 3.900 0.995 ;
        RECT  2.980 1.500 3.900 1.620 ;
        RECT  3.695 1.120 3.780 1.380 ;
        RECT  3.575 0.620 3.695 1.380 ;
        RECT  2.580 0.620 3.575 0.740 ;
        RECT  3.030 0.860 3.290 1.005 ;
        RECT  2.720 0.860 3.030 0.980 ;
        RECT  2.860 1.360 2.980 1.620 ;
        RECT  2.600 0.860 2.720 1.860 ;
        RECT  2.270 0.860 2.600 0.980 ;
        RECT  2.480 1.360 2.600 1.620 ;
        RECT  2.470 1.980 2.590 2.140 ;
        RECT  2.460 0.475 2.580 0.740 ;
        RECT  1.960 2.020 2.470 2.140 ;
        RECT  2.150 0.620 2.460 0.740 ;
        RECT  2.320 1.715 2.395 1.885 ;
        RECT  2.200 1.165 2.320 1.885 ;
        RECT  1.380 0.380 2.270 0.500 ;
        RECT  2.150 1.165 2.200 1.285 ;
        RECT  2.030 0.620 2.150 1.285 ;
        RECT  0.600 1.480 2.080 1.600 ;
        RECT  1.700 2.020 1.960 2.190 ;
        RECT  1.620 0.745 1.760 0.865 ;
        RECT  1.500 0.745 1.620 1.335 ;
        RECT  1.090 1.170 1.500 1.335 ;
        RECT  1.260 0.380 1.380 0.740 ;
        RECT  0.960 0.620 1.260 0.740 ;
        RECT  0.810 1.215 1.090 1.335 ;
        RECT  0.690 0.670 0.810 1.335 ;
        RECT  0.255 0.670 0.690 0.790 ;
        RECT  0.230 1.215 0.690 1.335 ;
        RECT  0.085 0.595 0.255 0.790 ;
        RECT  0.110 1.215 0.230 2.040 ;
    END
END EDFFX2AD
MACRO EDFFX4AD
    CLASS CORE ;
    FOREIGN EDFFX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.635 0.355 9.730 1.920 ;
        RECT  9.590 0.355 9.635 2.180 ;
        RECT  9.465 0.355 9.590 0.785 ;
        RECT  9.465 1.490 9.590 2.180 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.745 0.355 8.915 1.635 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.860 0.545 1.280 ;
        END
        AntennaGateArea 0.119 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.775 0.910 1.175 1.140 ;
        END
        AntennaGateArea 0.071 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.385 1.130 3.735 1.355 ;
        END
        AntennaGateArea 0.094 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.995 -0.210 10.080 0.210 ;
        RECT  9.850 -0.210 9.995 0.830 ;
        RECT  9.275 -0.210 9.850 0.210 ;
        RECT  9.105 -0.210 9.275 0.785 ;
        RECT  8.555 -0.210 9.105 0.210 ;
        RECT  8.385 -0.210 8.555 0.575 ;
        RECT  7.775 -0.210 8.385 0.210 ;
        RECT  7.515 -0.210 7.775 0.310 ;
        RECT  6.455 -0.210 7.515 0.210 ;
        RECT  6.195 -0.210 6.455 0.310 ;
        RECT  5.155 -0.210 6.195 0.210 ;
        RECT  4.895 -0.210 5.155 0.500 ;
        RECT  3.870 -0.210 4.895 0.210 ;
        RECT  3.350 -0.210 3.870 0.415 ;
        RECT  1.840 -0.210 3.350 0.210 ;
        RECT  1.580 -0.210 1.840 0.260 ;
        RECT  0.680 -0.210 1.580 0.210 ;
        RECT  0.420 -0.210 0.680 0.740 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.990 2.310 10.080 2.730 ;
        RECT  9.850 1.445 9.990 2.730 ;
        RECT  9.275 2.310 9.850 2.730 ;
        RECT  9.105 1.995 9.275 2.730 ;
        RECT  8.600 2.310 9.105 2.730 ;
        RECT  8.340 1.995 8.600 2.730 ;
        RECT  7.950 2.310 8.340 2.730 ;
        RECT  7.690 2.220 7.950 2.730 ;
        RECT  6.560 2.310 7.690 2.730 ;
        RECT  6.300 2.220 6.560 2.730 ;
        RECT  5.300 2.310 6.300 2.730 ;
        RECT  5.040 2.220 5.300 2.730 ;
        RECT  4.060 2.310 5.040 2.730 ;
        RECT  3.800 2.220 4.060 2.730 ;
        RECT  3.270 2.310 3.800 2.730 ;
        RECT  3.010 2.260 3.270 2.730 ;
        RECT  1.700 2.310 3.010 2.730 ;
        RECT  1.440 1.990 1.700 2.730 ;
        RECT  0.255 2.310 1.440 2.730 ;
        RECT  0.085 1.640 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.080 2.520 ;
        LAYER M1 ;
        RECT  9.260 1.020 9.460 1.280 ;
        RECT  9.140 1.020 9.260 1.875 ;
        RECT  8.625 1.755 9.140 1.875 ;
        RECT  8.505 0.695 8.625 1.875 ;
        RECT  8.125 0.695 8.505 0.815 ;
        RECT  8.130 1.400 8.505 1.520 ;
        RECT  7.650 1.080 8.385 1.210 ;
        RECT  8.010 1.400 8.130 2.100 ;
        RECT  7.955 0.525 8.125 0.815 ;
        RECT  2.900 1.980 8.010 2.100 ;
        RECT  7.530 0.430 7.650 1.850 ;
        RECT  5.805 0.430 7.530 0.550 ;
        RECT  5.670 1.730 7.530 1.850 ;
        RECT  7.290 0.670 7.410 1.610 ;
        RECT  6.865 0.670 7.290 0.790 ;
        RECT  7.050 0.910 7.170 1.560 ;
        RECT  5.945 1.440 7.050 1.560 ;
        RECT  6.745 0.670 6.865 1.315 ;
        RECT  6.205 1.195 6.745 1.315 ;
        RECT  6.445 0.950 6.585 1.070 ;
        RECT  6.325 0.670 6.445 1.070 ;
        RECT  5.325 0.670 6.325 0.790 ;
        RECT  6.085 0.910 6.205 1.315 ;
        RECT  5.565 0.910 6.085 1.030 ;
        RECT  5.815 1.200 5.945 1.610 ;
        RECT  5.295 1.490 5.815 1.610 ;
        RECT  5.545 0.380 5.805 0.550 ;
        RECT  5.445 0.910 5.565 1.370 ;
        RECT  4.890 1.250 5.445 1.370 ;
        RECT  5.065 0.620 5.325 1.105 ;
        RECT  5.175 1.490 5.295 1.860 ;
        RECT  2.970 1.740 5.175 1.860 ;
        RECT  4.305 0.620 5.065 0.740 ;
        RECT  4.630 1.250 4.890 1.620 ;
        RECT  4.545 0.860 4.775 0.980 ;
        RECT  4.545 1.250 4.630 1.370 ;
        RECT  4.425 0.860 4.545 1.370 ;
        RECT  4.305 1.500 4.370 1.620 ;
        RECT  4.185 0.620 4.305 1.620 ;
        RECT  4.095 0.620 4.185 1.000 ;
        RECT  3.220 1.500 4.185 1.620 ;
        RECT  3.975 1.120 4.065 1.380 ;
        RECT  3.855 0.545 3.975 1.380 ;
        RECT  2.860 0.545 3.855 0.665 ;
        RECT  2.970 0.860 3.560 1.005 ;
        RECT  3.100 1.360 3.220 1.620 ;
        RECT  2.850 0.860 2.970 1.860 ;
        RECT  2.780 1.980 2.900 2.140 ;
        RECT  2.740 0.460 2.860 0.740 ;
        RECT  2.550 0.860 2.850 1.005 ;
        RECT  2.690 1.360 2.850 1.620 ;
        RECT  2.180 2.020 2.780 2.140 ;
        RECT  2.425 0.620 2.740 0.740 ;
        RECT  2.515 1.750 2.730 1.870 ;
        RECT  1.690 0.380 2.550 0.500 ;
        RECT  2.425 1.160 2.515 1.870 ;
        RECT  2.395 0.620 2.425 1.870 ;
        RECT  2.305 0.620 2.395 1.280 ;
        RECT  2.155 1.610 2.275 1.870 ;
        RECT  1.920 2.020 2.180 2.190 ;
        RECT  0.930 1.750 2.155 1.870 ;
        RECT  1.930 0.840 2.070 0.960 ;
        RECT  1.810 0.840 1.930 1.125 ;
        RECT  1.460 1.005 1.810 1.125 ;
        RECT  1.570 0.380 1.690 0.740 ;
        RECT  1.030 0.620 1.570 0.740 ;
        RECT  1.340 1.005 1.460 1.520 ;
        RECT  0.225 1.400 1.340 1.520 ;
        RECT  0.760 1.750 0.930 1.945 ;
        RECT  0.225 0.595 0.275 0.765 ;
        RECT  0.105 0.595 0.225 1.520 ;
    END
END EDFFX4AD
MACRO EDFFXLAD
    CLASS CORE ;
    FOREIGN EDFFXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 1.425 7.490 1.685 ;
        RECT  7.330 0.555 7.450 1.685 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.850 0.865 6.970 1.860 ;
        RECT  6.730 0.865 6.850 1.095 ;
        RECT  6.260 1.740 6.850 1.860 ;
        RECT  6.610 0.555 6.730 1.095 ;
        END
        AntennaDiffArea 0.134 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.170 0.910 0.570 1.095 ;
        END
        AntennaGateArea 0.119 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.930 0.865 1.375 1.050 ;
        END
        AntennaGateArea 0.071 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.100 1.130 3.455 1.355 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.160 -0.210 7.560 0.210 ;
        RECT  6.900 -0.210 7.160 0.745 ;
        RECT  6.140 -0.210 6.900 0.210 ;
        RECT  5.880 -0.210 6.140 0.445 ;
        RECT  4.685 -0.210 5.880 0.210 ;
        RECT  4.425 -0.210 4.685 0.415 ;
        RECT  3.470 -0.210 4.425 0.210 ;
        RECT  3.210 -0.210 3.470 0.415 ;
        RECT  1.575 -0.210 3.210 0.210 ;
        RECT  1.405 -0.210 1.575 0.260 ;
        RECT  0.545 -0.210 1.405 0.210 ;
        RECT  0.375 -0.210 0.545 0.335 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.140 2.310 7.560 2.730 ;
        RECT  6.880 2.220 7.140 2.730 ;
        RECT  6.140 2.310 6.880 2.730 ;
        RECT  5.880 2.220 6.140 2.730 ;
        RECT  4.890 2.310 5.880 2.730 ;
        RECT  4.630 2.220 4.890 2.730 ;
        RECT  3.780 2.310 4.630 2.730 ;
        RECT  3.520 2.220 3.780 2.730 ;
        RECT  3.060 2.310 3.520 2.730 ;
        RECT  2.800 2.250 3.060 2.730 ;
        RECT  1.425 2.310 2.800 2.730 ;
        RECT  1.255 1.720 1.425 2.730 ;
        RECT  0.610 2.310 1.255 2.730 ;
        RECT  0.490 2.055 0.610 2.730 ;
        RECT  0.000 2.310 0.490 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  7.090 1.005 7.210 2.100 ;
        RECT  5.900 1.980 7.090 2.100 ;
        RECT  6.610 1.330 6.730 1.590 ;
        RECT  6.490 1.330 6.610 1.450 ;
        RECT  6.370 0.755 6.490 1.450 ;
        RECT  6.170 0.755 6.370 0.875 ;
        RECT  5.900 1.330 6.370 1.450 ;
        RECT  6.080 1.000 6.250 1.210 ;
        RECT  5.640 1.000 6.080 1.120 ;
        RECT  5.780 1.300 5.900 2.100 ;
        RECT  2.590 1.980 5.780 2.100 ;
        RECT  5.520 0.755 5.640 1.800 ;
        RECT  5.360 0.375 5.620 0.570 ;
        RECT  5.290 0.755 5.520 1.015 ;
        RECT  5.260 1.680 5.520 1.800 ;
        RECT  5.170 1.385 5.400 1.520 ;
        RECT  5.170 0.450 5.360 0.570 ;
        RECT  5.050 0.450 5.170 1.520 ;
        RECT  4.750 1.085 5.050 1.205 ;
        RECT  4.805 0.395 4.925 0.655 ;
        RECT  4.020 0.535 4.805 0.655 ;
        RECT  4.630 1.085 4.750 1.860 ;
        RECT  4.510 1.085 4.630 1.345 ;
        RECT  2.720 1.740 4.630 1.860 ;
        RECT  4.380 1.500 4.510 1.620 ;
        RECT  4.250 0.810 4.380 1.620 ;
        RECT  4.210 0.810 4.250 1.320 ;
        RECT  4.140 1.060 4.210 1.320 ;
        RECT  4.020 1.500 4.130 1.620 ;
        RECT  3.900 0.535 4.020 1.620 ;
        RECT  3.815 0.535 3.900 0.995 ;
        RECT  2.980 1.500 3.900 1.620 ;
        RECT  3.695 1.120 3.780 1.380 ;
        RECT  3.575 0.620 3.695 1.380 ;
        RECT  2.580 0.620 3.575 0.740 ;
        RECT  3.030 0.860 3.290 1.005 ;
        RECT  2.720 0.860 3.030 0.980 ;
        RECT  2.860 1.360 2.980 1.620 ;
        RECT  2.600 0.860 2.720 1.860 ;
        RECT  2.270 0.860 2.600 0.980 ;
        RECT  2.480 1.360 2.600 1.620 ;
        RECT  2.470 1.980 2.590 2.140 ;
        RECT  2.460 0.475 2.580 0.740 ;
        RECT  1.960 2.020 2.470 2.140 ;
        RECT  2.150 0.620 2.460 0.740 ;
        RECT  2.320 1.715 2.395 1.885 ;
        RECT  2.200 1.165 2.320 1.885 ;
        RECT  1.380 0.380 2.270 0.500 ;
        RECT  2.150 1.165 2.200 1.285 ;
        RECT  2.030 0.620 2.150 1.285 ;
        RECT  0.600 1.480 2.080 1.600 ;
        RECT  1.700 2.020 1.960 2.190 ;
        RECT  1.620 0.745 1.760 0.865 ;
        RECT  1.500 0.745 1.620 1.335 ;
        RECT  1.090 1.170 1.500 1.335 ;
        RECT  1.260 0.380 1.380 0.740 ;
        RECT  0.960 0.620 1.260 0.740 ;
        RECT  0.810 1.215 1.090 1.335 ;
        RECT  0.690 0.670 0.810 1.335 ;
        RECT  0.255 0.670 0.690 0.790 ;
        RECT  0.230 1.215 0.690 1.335 ;
        RECT  0.085 0.595 0.255 0.790 ;
        RECT  0.110 1.215 0.230 2.040 ;
    END
END EDFFXLAD
MACRO FILL16AD
    CLASS CORE SPACER ;
    FOREIGN FILL16AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.595 -0.210 4.480 0.210 ;
        RECT  3.595 0.445 3.960 0.615 ;
        RECT  3.075 -0.210 3.595 0.615 ;
        RECT  1.380 -0.210 3.075 0.210 ;
        RECT  2.710 0.445 3.075 0.615 ;
        RECT  1.380 0.445 1.745 0.615 ;
        RECT  0.860 -0.210 1.380 0.615 ;
        RECT  0.000 -0.210 0.860 0.210 ;
        RECT  0.495 0.445 0.860 0.615 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.555 2.310 4.480 2.730 ;
        RECT  3.555 1.900 3.920 2.070 ;
        RECT  3.035 1.900 3.555 2.730 ;
        RECT  2.670 1.900 3.035 2.070 ;
        RECT  1.455 2.310 3.035 2.730 ;
        RECT  1.455 1.900 1.820 2.070 ;
        RECT  0.935 1.900 1.455 2.730 ;
        RECT  0.570 1.900 0.935 2.070 ;
        RECT  0.000 2.310 0.935 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
	 END
END FILL16AD
MACRO FILL1AD
    CLASS CORE SPACER ;
    FOREIGN FILL1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.280 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.210 0.280 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.310 0.280 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 0.280 2.520 ;
	 END
END FILL1AD
MACRO FILL2AD
    CLASS CORE SPACER ;
    FOREIGN FILL2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.410 -0.210 0.560 0.210 ;
        RECT  0.150 -0.210 0.410 0.590 ;
        RECT  0.000 -0.210 0.150 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.410 2.310 0.560 2.730 ;
        RECT  0.150 1.930 0.410 2.730 ;
        RECT  0.000 2.310 0.150 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 0.560 2.520 ;
	 END
END FILL2AD
MACRO FILL32AD
    CLASS CORE SPACER ;
    FOREIGN FILL32AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.020 -0.210 8.960 0.210 ;
        RECT  8.020 0.445 8.410 0.615 ;
        RECT  7.555 -0.210 8.020 0.615 ;
        RECT  5.795 -0.210 7.555 0.210 ;
        RECT  7.160 0.445 7.555 0.615 ;
        RECT  5.795 0.445 6.195 0.615 ;
        RECT  5.330 -0.210 5.795 0.615 ;
        RECT  3.565 -0.210 5.330 0.210 ;
        RECT  4.945 0.445 5.330 0.615 ;
        RECT  3.565 0.445 3.960 0.615 ;
        RECT  3.100 -0.210 3.565 0.615 ;
        RECT  1.355 -0.210 3.100 0.210 ;
        RECT  2.710 0.445 3.100 0.615 ;
        RECT  1.355 0.445 1.745 0.615 ;
        RECT  0.890 -0.210 1.355 0.615 ;
        RECT  0.000 -0.210 0.890 0.210 ;
        RECT  0.495 0.445 0.890 0.615 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.980 2.310 8.960 2.730 ;
        RECT  7.980 1.905 8.370 2.075 ;
        RECT  7.515 1.905 7.980 2.730 ;
        RECT  7.120 1.905 7.515 2.075 ;
        RECT  5.875 2.310 7.515 2.730 ;
        RECT  5.875 1.905 6.270 2.075 ;
        RECT  5.410 1.905 5.875 2.730 ;
        RECT  5.020 1.905 5.410 2.075 ;
        RECT  3.525 2.310 5.410 2.730 ;
        RECT  3.525 1.905 3.920 2.075 ;
        RECT  3.060 1.905 3.525 2.730 ;
        RECT  2.670 1.905 3.060 2.075 ;
        RECT  1.435 2.310 3.060 2.730 ;
        RECT  1.435 1.905 1.820 2.075 ;
        RECT  0.970 1.905 1.435 2.730 ;
        RECT  0.570 1.905 0.970 2.075 ;
        RECT  0.000 2.310 0.970 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.960 2.520 ;
	 END
END FILL32AD
MACRO FILL4AD
    CLASS CORE SPACER ;
    FOREIGN FILL4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.640 -0.210 1.120 0.210 ;
        RECT  0.470 -0.210 0.640 0.615 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.620 2.310 1.120 2.730 ;
        RECT  0.450 1.905 0.620 2.730 ;
        RECT  0.000 2.310 0.450 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
	 END
END FILL4AD
MACRO FILL64AD
    CLASS CORE SPACER ;
    FOREIGN FILL64AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.960 -0.210 17.920 0.210 ;
        RECT  16.960 0.445 17.265 0.615 ;
        RECT  16.540 -0.210 16.960 0.615 ;
        RECT  14.860 -0.210 16.540 0.210 ;
        RECT  16.315 0.445 16.540 0.615 ;
        RECT  14.860 0.445 15.050 0.615 ;
        RECT  14.440 -0.210 14.860 0.615 ;
        RECT  12.510 -0.210 14.440 0.210 ;
        RECT  14.100 0.445 14.440 0.615 ;
        RECT  12.510 0.445 12.815 0.615 ;
        RECT  12.090 -0.210 12.510 0.615 ;
        RECT  10.410 -0.210 12.090 0.210 ;
        RECT  11.865 0.445 12.090 0.615 ;
        RECT  10.410 0.445 10.600 0.615 ;
        RECT  9.990 -0.210 10.410 0.615 ;
        RECT  7.955 -0.210 9.990 0.210 ;
        RECT  9.650 0.445 9.990 0.615 ;
        RECT  7.955 0.445 8.260 0.615 ;
        RECT  7.535 -0.210 7.955 0.615 ;
        RECT  5.855 -0.210 7.535 0.210 ;
        RECT  7.310 0.445 7.535 0.615 ;
        RECT  5.855 0.445 6.045 0.615 ;
        RECT  5.435 -0.210 5.855 0.615 ;
        RECT  3.505 -0.210 5.435 0.210 ;
        RECT  5.095 0.445 5.435 0.615 ;
        RECT  3.505 0.470 3.855 0.590 ;
        RECT  3.085 -0.210 3.505 0.590 ;
        RECT  1.405 -0.210 3.085 0.210 ;
        RECT  2.815 0.470 3.085 0.590 ;
        RECT  1.405 0.445 1.595 0.615 ;
        RECT  0.985 -0.210 1.405 0.615 ;
        RECT  0.000 -0.210 0.985 0.210 ;
        RECT  0.645 0.445 0.985 0.615 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.960 2.310 17.920 2.730 ;
        RECT  16.960 1.905 17.225 2.075 ;
        RECT  16.540 1.905 16.960 2.730 ;
        RECT  16.275 1.905 16.540 2.075 ;
        RECT  14.860 2.310 16.540 2.730 ;
        RECT  14.860 1.905 15.125 2.075 ;
        RECT  14.440 1.905 14.860 2.730 ;
        RECT  14.175 1.905 14.440 2.075 ;
        RECT  12.510 2.310 14.440 2.730 ;
        RECT  12.510 1.905 12.775 2.075 ;
        RECT  12.090 1.905 12.510 2.730 ;
        RECT  11.825 1.905 12.090 2.075 ;
        RECT  10.410 2.310 12.090 2.730 ;
        RECT  10.410 1.905 10.675 2.075 ;
        RECT  9.990 1.905 10.410 2.730 ;
        RECT  9.725 1.905 9.990 2.075 ;
        RECT  7.955 2.310 9.990 2.730 ;
        RECT  7.955 1.905 8.220 2.075 ;
        RECT  7.535 1.905 7.955 2.730 ;
        RECT  7.270 1.905 7.535 2.075 ;
        RECT  5.855 2.310 7.535 2.730 ;
        RECT  5.855 1.905 6.120 2.075 ;
        RECT  5.435 1.905 5.855 2.730 ;
        RECT  5.170 1.905 5.435 2.075 ;
        RECT  3.505 2.310 5.435 2.730 ;
        RECT  3.505 1.905 3.770 2.075 ;
        RECT  3.085 1.905 3.505 2.730 ;
        RECT  2.820 1.905 3.085 2.075 ;
        RECT  1.405 2.310 3.085 2.730 ;
        RECT  1.405 1.905 1.670 2.075 ;
        RECT  0.985 1.905 1.405 2.730 ;
        RECT  0.720 1.905 0.985 2.075 ;
        RECT  0.000 2.310 0.985 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 17.920 2.520 ;
	 END
END FILL64AD
MACRO FILL8AD
    CLASS CORE SPACER ;
    FOREIGN FILL8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.390 -0.210 2.240 0.210 ;
        RECT  1.390 0.445 1.745 0.615 ;
        RECT  0.870 -0.210 1.390 0.620 ;
        RECT  0.000 -0.210 0.870 0.210 ;
        RECT  0.495 0.445 0.870 0.615 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.390 2.310 2.240 2.730 ;
        RECT  1.390 1.900 1.755 2.070 ;
        RECT  0.870 1.900 1.390 2.730 ;
        RECT  0.505 1.900 0.870 2.070 ;
        RECT  0.000 2.310 0.870 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
	 END
END FILL8AD
MACRO FILLCAP16AD
    CLASS CORE SPACER ;
    FOREIGN FILLCAP16AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.045 -0.210 4.200 0.210 ;
        RECT  3.875 -0.210 4.045 0.795 ;
        RECT  0.425 -0.210 3.875 0.210 ;
        RECT  0.255 -0.210 0.425 0.805 ;
        RECT  0.000 -0.210 0.255 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.045 2.310 4.200 2.730 ;
        RECT  3.875 1.660 4.045 2.730 ;
        RECT  0.425 2.310 3.875 2.730 ;
        RECT  0.255 1.735 0.425 2.730 ;
        RECT  0.000 2.310 0.255 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  3.245 0.890 3.765 1.550 ;
        RECT  2.235 1.430 3.245 1.550 ;
        RECT  2.210 1.190 2.790 1.310 ;
        RECT  2.210 0.365 2.235 0.795 ;
        RECT  2.065 1.430 2.235 1.945 ;
        RECT  2.090 0.365 2.210 1.310 ;
        RECT  2.065 0.365 2.090 0.795 ;
        RECT  1.510 1.190 2.090 1.310 ;
        RECT  1.055 1.430 2.065 1.550 ;
        RECT  0.535 0.890 1.055 1.550 ;
    END
END FILLCAP16AD
MACRO FILLCAP32AD
    CLASS CORE SPACER ;
    FOREIGN FILLCAP32AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.905 -0.210 8.120 0.210 ;
        RECT  7.735 -0.210 7.905 0.785 ;
        RECT  4.160 -0.210 7.735 0.210 ;
        RECT  3.900 -0.210 4.160 0.500 ;
        RECT  0.325 -0.210 3.900 0.210 ;
        RECT  0.155 -0.210 0.325 0.785 ;
        RECT  0.000 -0.210 0.155 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.905 2.310 8.120 2.730 ;
        RECT  7.735 1.735 7.905 2.730 ;
        RECT  4.115 2.310 7.735 2.730 ;
        RECT  3.945 1.735 4.115 2.730 ;
        RECT  0.325 2.310 3.945 2.730 ;
        RECT  0.155 1.535 0.325 2.730 ;
        RECT  0.000 2.310 0.155 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.120 2.520 ;
        LAYER M1 ;
        RECT  7.105 0.890 7.625 1.550 ;
        RECT  6.015 1.430 7.105 1.550 ;
        RECT  6.015 1.190 6.830 1.310 ;
        RECT  5.845 0.370 6.015 1.310 ;
        RECT  5.845 1.430 6.015 1.975 ;
        RECT  2.215 0.620 5.845 0.740 ;
        RECT  5.290 1.190 5.845 1.310 ;
        RECT  4.930 1.430 5.845 1.550 ;
        RECT  3.130 0.920 4.930 1.550 ;
        RECT  2.215 1.430 3.130 1.550 ;
        RECT  2.215 1.190 2.770 1.310 ;
        RECT  2.045 0.365 2.215 1.310 ;
        RECT  2.045 1.430 2.215 1.945 ;
        RECT  1.230 1.190 2.045 1.310 ;
        RECT  1.005 1.430 2.045 1.550 ;
        RECT  0.485 0.900 1.005 1.550 ;
    END
END FILLCAP32AD
MACRO FILLCAP3AD
    CLASS CORE SPACER ;
    FOREIGN FILLCAP3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.285 -0.210 0.840 0.210 ;
        RECT  0.115 -0.210 0.285 0.655 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.725 2.310 0.840 2.730 ;
        RECT  0.555 1.585 0.725 2.730 ;
        RECT  0.000 2.310 0.555 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 0.840 2.520 ;
        LAYER M1 ;
        RECT  0.610 0.485 0.730 1.325 ;
        RECT  0.555 0.485 0.610 0.655 ;
        RECT  0.360 1.205 0.610 1.325 ;
        RECT  0.235 0.900 0.490 1.020 ;
        RECT  0.235 1.585 0.285 2.015 ;
        RECT  0.115 0.900 0.235 2.015 ;
    END
END FILLCAP3AD
MACRO FILLCAP4AD
    CLASS CORE SPACER ;
    FOREIGN FILLCAP4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.285 -0.210 1.120 0.210 ;
        RECT  0.115 -0.210 0.285 0.825 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.005 2.310 1.120 2.730 ;
        RECT  0.835 1.530 1.005 2.730 ;
        RECT  0.000 2.310 0.835 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
        LAYER M1 ;
        RECT  0.955 0.400 1.005 0.830 ;
        RECT  0.835 0.400 0.955 1.330 ;
        RECT  0.610 1.210 0.835 1.330 ;
        RECT  0.235 0.950 0.540 1.070 ;
        RECT  0.235 1.545 0.285 1.975 ;
        RECT  0.115 0.950 0.235 1.975 ;
    END
END FILLCAP4AD
MACRO FILLCAP64AD
    CLASS CORE SPACER ;
    FOREIGN FILLCAP64AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  17.105 -0.210 17.360 0.210 ;
        RECT  16.935 -0.210 17.105 0.575 ;
        RECT  13.070 -0.210 16.935 0.210 ;
        RECT  13.070 0.380 13.100 0.500 ;
        RECT  12.870 -0.210 13.070 0.500 ;
        RECT  8.730 -0.210 12.870 0.210 ;
        RECT  12.840 0.380 12.870 0.500 ;
        RECT  8.730 0.375 8.845 0.545 ;
        RECT  8.530 -0.210 8.730 0.545 ;
        RECT  4.420 -0.210 8.530 0.210 ;
        RECT  8.415 0.375 8.530 0.545 ;
        RECT  4.160 -0.210 4.420 0.500 ;
        RECT  0.325 -0.210 4.160 0.210 ;
        RECT  0.155 -0.210 0.325 0.710 ;
        RECT  0.000 -0.210 0.155 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  17.105 2.310 17.360 2.730 ;
        RECT  16.935 1.670 17.105 2.730 ;
        RECT  13.055 2.310 16.935 2.730 ;
        RECT  12.885 1.735 13.055 2.730 ;
        RECT  8.840 2.310 12.885 2.730 ;
        RECT  8.840 1.620 8.975 2.150 ;
        RECT  8.420 1.620 8.840 2.730 ;
        RECT  8.285 1.620 8.420 2.150 ;
        RECT  4.375 2.310 8.420 2.730 ;
        RECT  4.205 1.735 4.375 2.730 ;
        RECT  0.325 2.310 4.205 2.730 ;
        RECT  0.155 1.665 0.325 2.730 ;
        RECT  0.000 2.310 0.155 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 17.360 2.520 ;
        LAYER M1 ;
        RECT  16.910 1.430 17.130 1.550 ;
        RECT  16.130 0.920 16.910 1.550 ;
        RECT  15.085 1.430 16.130 1.550 ;
        RECT  15.085 1.190 15.640 1.310 ;
        RECT  14.915 0.355 15.085 1.310 ;
        RECT  14.915 1.430 15.085 1.960 ;
        RECT  11.025 0.620 14.915 0.740 ;
        RECT  14.360 1.190 14.915 1.310 ;
        RECT  13.870 1.430 14.915 1.550 ;
        RECT  12.330 0.920 13.870 1.550 ;
        RECT  11.025 1.430 12.330 1.550 ;
        RECT  11.000 1.190 11.840 1.310 ;
        RECT  11.000 0.365 11.025 0.795 ;
        RECT  10.855 1.430 11.025 1.945 ;
        RECT  10.880 0.365 11.000 1.310 ;
        RECT  10.855 0.365 10.880 0.795 ;
        RECT  10.300 1.190 10.880 1.310 ;
        RECT  9.130 0.620 10.855 0.740 ;
        RECT  9.770 1.430 10.855 1.550 ;
        RECT  9.250 0.920 9.770 1.550 ;
        RECT  8.010 1.320 9.250 1.440 ;
        RECT  9.010 0.620 9.130 0.810 ;
        RECT  8.250 0.690 9.010 0.810 ;
        RECT  8.130 0.620 8.250 0.810 ;
        RECT  6.405 0.620 8.130 0.740 ;
        RECT  7.490 0.920 8.010 1.550 ;
        RECT  6.405 1.430 7.490 1.550 ;
        RECT  6.380 1.190 7.220 1.310 ;
        RECT  6.380 0.375 6.405 0.805 ;
        RECT  6.235 1.430 6.405 1.945 ;
        RECT  6.260 0.375 6.380 1.310 ;
        RECT  6.235 0.375 6.260 0.805 ;
        RECT  5.680 1.190 6.260 1.310 ;
        RECT  2.345 0.620 6.235 0.740 ;
        RECT  5.190 1.430 6.235 1.550 ;
        RECT  3.650 0.920 5.190 1.550 ;
        RECT  2.345 1.430 3.650 1.550 ;
        RECT  2.345 1.190 3.160 1.310 ;
        RECT  2.175 0.375 2.345 1.310 ;
        RECT  2.175 1.430 2.345 1.945 ;
        RECT  1.620 1.190 2.175 1.310 ;
        RECT  1.215 1.430 2.175 1.550 ;
        RECT  0.435 0.920 1.215 1.550 ;
    END
END FILLCAP64AD
MACRO FILLCAP8AD
    CLASS CORE SPACER ;
    FOREIGN FILLCAP8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.325 -0.210 1.960 0.210 ;
        RECT  0.155 -0.210 0.325 0.785 ;
        RECT  0.000 -0.210 0.155 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.815 2.310 1.960 2.730 ;
        RECT  1.645 1.565 1.815 2.730 ;
        RECT  0.000 2.310 1.645 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.775 0.375 1.825 0.805 ;
        RECT  1.655 0.375 1.775 1.305 ;
        RECT  1.100 1.185 1.655 1.305 ;
        RECT  0.325 0.925 0.870 1.045 ;
        RECT  0.205 0.925 0.325 1.995 ;
        RECT  0.155 1.565 0.205 1.995 ;
    END
END FILLCAP8AD
MACRO INVX10AD
    CLASS CORE ;
    FOREIGN INVX10AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.930 0.390 2.130 0.895 ;
        RECT  1.945 1.375 2.115 2.090 ;
        RECT  1.785 1.375 1.945 1.665 ;
        RECT  1.785 0.630 1.930 0.895 ;
        RECT  1.390 0.630 1.785 1.665 ;
        RECT  1.365 0.630 1.390 2.080 ;
        RECT  1.260 0.390 1.365 2.080 ;
        RECT  1.195 0.390 1.260 0.895 ;
        RECT  1.170 1.375 1.260 2.080 ;
        RECT  0.645 0.615 1.195 0.895 ;
        RECT  0.670 1.375 1.170 1.665 ;
        RECT  0.450 1.375 0.670 2.080 ;
        RECT  0.475 0.390 0.645 0.895 ;
        END
        AntennaDiffArea 1.217 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.065 1.090 1.185 ;
        RECT  0.070 0.865 0.210 1.185 ;
        END
        AntennaGateArea 0.81 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.210 2.240 0.210 ;
        RECT  1.555 -0.210 1.725 0.495 ;
        RECT  1.005 -0.210 1.555 0.210 ;
        RECT  0.835 -0.210 1.005 0.495 ;
        RECT  0.290 -0.210 0.835 0.210 ;
        RECT  0.110 -0.210 0.290 0.730 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.760 2.310 2.240 2.730 ;
        RECT  1.540 1.845 1.760 2.730 ;
        RECT  1.030 2.310 1.540 2.730 ;
        RECT  0.810 1.845 1.030 2.730 ;
        RECT  0.285 2.310 0.810 2.730 ;
        RECT  0.115 1.585 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
	 END
END INVX10AD
MACRO INVX12AD
    CLASS CORE ;
    FOREIGN INVX12AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.905 0.420 2.075 2.110 ;
        RECT  1.880 0.655 1.905 2.110 ;
        RECT  1.360 0.655 1.880 1.630 ;
        RECT  1.140 0.395 1.360 2.110 ;
        RECT  1.125 0.670 1.140 1.675 ;
        RECT  0.640 0.670 1.125 0.895 ;
        RECT  0.640 1.405 1.125 1.675 ;
        RECT  0.420 0.420 0.640 0.895 ;
        RECT  0.420 1.405 0.640 2.110 ;
        END
        AntennaDiffArea 1.266 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.065 0.990 1.230 ;
        RECT  0.070 1.065 0.210 1.375 ;
        END
        AntennaGateArea 0.972 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 -0.210 2.520 0.210 ;
        RECT  2.265 -0.210 2.435 0.910 ;
        RECT  1.760 -0.210 2.265 0.210 ;
        RECT  1.500 -0.210 1.760 0.525 ;
        RECT  1.020 -0.210 1.500 0.210 ;
        RECT  0.760 -0.210 1.020 0.525 ;
        RECT  0.255 -0.210 0.760 0.210 ;
        RECT  0.085 -0.210 0.255 0.865 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 2.310 2.520 2.730 ;
        RECT  2.265 1.420 2.435 2.730 ;
        RECT  1.740 2.310 2.265 2.730 ;
        RECT  1.480 1.760 1.740 2.730 ;
        RECT  1.020 2.310 1.480 2.730 ;
        RECT  0.760 1.855 1.020 2.730 ;
        RECT  0.255 2.310 0.760 2.730 ;
        RECT  0.085 1.680 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
	 END
END INVX12AD
MACRO INVX14AD
    CLASS CORE ;
    FOREIGN INVX14AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.745 0.360 2.915 2.065 ;
        RECT  2.190 0.890 2.745 1.665 ;
        RECT  2.165 0.385 2.190 1.665 ;
        RECT  1.995 0.385 2.165 2.065 ;
        RECT  1.970 0.385 1.995 1.665 ;
        RECT  1.430 0.640 1.970 1.665 ;
        RECT  1.210 0.385 1.430 0.890 ;
        RECT  1.405 1.375 1.430 1.665 ;
        RECT  1.235 1.375 1.405 2.065 ;
        RECT  0.645 1.375 1.235 1.665 ;
        RECT  0.670 0.615 1.210 0.890 ;
        RECT  0.450 0.360 0.670 0.890 ;
        RECT  0.475 1.375 0.645 2.065 ;
        END
        AntennaDiffArea 1.735 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 1.070 1.310 1.190 ;
        RECT  0.070 0.860 0.230 1.190 ;
        END
        AntennaGateArea 1.134 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.570 -0.210 3.080 0.210 ;
        RECT  2.350 -0.210 2.570 0.675 ;
        RECT  1.830 -0.210 2.350 0.210 ;
        RECT  1.570 -0.210 1.830 0.510 ;
        RECT  1.070 -0.210 1.570 0.210 ;
        RECT  0.810 -0.210 1.070 0.495 ;
        RECT  0.290 -0.210 0.810 0.210 ;
        RECT  0.105 -0.210 0.290 0.700 ;
        RECT  0.000 -0.210 0.105 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.570 2.310 3.080 2.730 ;
        RECT  2.350 1.845 2.570 2.730 ;
        RECT  1.810 2.310 2.350 2.730 ;
        RECT  1.590 1.845 1.810 2.730 ;
        RECT  1.050 2.310 1.590 2.730 ;
        RECT  0.830 1.845 1.050 2.730 ;
        RECT  0.275 2.310 0.830 2.730 ;
        RECT  0.100 1.370 0.275 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
	 END
END INVX14AD
MACRO INVX16AD
    CLASS CORE ;
    FOREIGN INVX16AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.610 0.400 2.830 2.065 ;
        RECT  2.110 0.830 2.610 1.630 ;
        RECT  2.105 0.400 2.110 1.630 ;
        RECT  1.890 0.400 2.105 2.065 ;
        RECT  1.410 0.830 1.890 1.630 ;
        RECT  1.390 0.375 1.410 1.630 ;
        RECT  1.220 0.375 1.390 2.065 ;
        RECT  1.170 0.375 1.220 0.890 ;
        RECT  1.170 1.375 1.220 2.065 ;
        RECT  0.670 0.630 1.170 0.890 ;
        RECT  0.645 1.375 1.170 1.625 ;
        RECT  0.450 0.375 0.670 0.890 ;
        RECT  0.475 1.375 0.645 2.065 ;
        END
        AntennaDiffArea 1.736 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.075 1.060 1.195 ;
        RECT  0.070 0.865 0.210 1.195 ;
        END
        AntennaGateArea 1.296 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.195 -0.210 3.360 0.210 ;
        RECT  3.025 -0.210 3.195 0.695 ;
        RECT  2.470 -0.210 3.025 0.210 ;
        RECT  2.250 -0.210 2.470 0.675 ;
        RECT  1.750 -0.210 2.250 0.210 ;
        RECT  1.530 -0.210 1.750 0.675 ;
        RECT  1.050 -0.210 1.530 0.210 ;
        RECT  0.790 -0.210 1.050 0.510 ;
        RECT  0.285 -0.210 0.790 0.210 ;
        RECT  0.115 -0.210 0.285 0.740 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.195 2.310 3.360 2.730 ;
        RECT  3.025 1.450 3.195 2.730 ;
        RECT  2.470 2.310 3.025 2.730 ;
        RECT  2.250 1.785 2.470 2.730 ;
        RECT  1.750 2.310 2.250 2.730 ;
        RECT  1.530 1.785 1.750 2.730 ;
        RECT  1.030 2.310 1.530 2.730 ;
        RECT  0.810 1.785 1.030 2.730 ;
        RECT  0.285 2.310 0.810 2.730 ;
        RECT  0.115 1.450 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
	 END
END INVX16AD
MACRO INVX18AD
    CLASS CORE ;
    FOREIGN INVX18AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.335 0.400 3.540 2.120 ;
        RECT  2.815 0.890 3.335 1.630 ;
        RECT  2.790 0.400 2.815 1.630 ;
        RECT  2.590 0.400 2.790 2.120 ;
        RECT  2.075 0.890 2.590 1.630 ;
        RECT  1.860 0.400 2.075 2.120 ;
        RECT  1.615 0.630 1.860 1.630 ;
        RECT  1.360 0.630 1.615 0.890 ;
        RECT  1.360 1.370 1.615 1.630 ;
        RECT  1.140 0.375 1.360 0.890 ;
        RECT  1.140 1.370 1.360 2.145 ;
        RECT  0.640 0.630 1.140 0.890 ;
        RECT  0.640 1.370 1.140 1.640 ;
        RECT  0.420 0.375 0.640 0.890 ;
        RECT  0.430 1.370 0.640 2.145 ;
        END
        AntennaDiffArea 2.109 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 1.070 1.455 1.190 ;
        RECT  0.070 0.860 0.230 1.190 ;
        END
        AntennaGateArea 1.458 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.190 -0.210 3.640 0.210 ;
        RECT  2.970 -0.210 3.190 0.675 ;
        RECT  2.440 -0.210 2.970 0.210 ;
        RECT  2.220 -0.210 2.440 0.675 ;
        RECT  1.740 -0.210 2.220 0.210 ;
        RECT  1.480 -0.210 1.740 0.485 ;
        RECT  1.020 -0.210 1.480 0.210 ;
        RECT  0.760 -0.210 1.020 0.485 ;
        RECT  0.255 -0.210 0.760 0.210 ;
        RECT  0.085 -0.210 0.255 0.700 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.190 2.310 3.640 2.730 ;
        RECT  2.970 1.760 3.190 2.730 ;
        RECT  2.445 2.310 2.970 2.730 ;
        RECT  2.225 1.760 2.445 2.730 ;
        RECT  1.720 2.310 2.225 2.730 ;
        RECT  1.500 1.760 1.720 2.730 ;
        RECT  1.000 2.310 1.500 2.730 ;
        RECT  0.780 1.760 1.000 2.730 ;
        RECT  0.255 2.310 0.780 2.730 ;
        RECT  0.085 1.405 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
	 END
END INVX18AD
MACRO INVX1AD
    CLASS CORE ;
    FOREIGN INVX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.675 0.640 0.770 1.525 ;
        RECT  0.610 0.640 0.675 1.925 ;
        RECT  0.535 0.640 0.610 0.900 ;
        RECT  0.515 1.365 0.610 1.925 ;
        END
        AntennaDiffArea 0.215 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.050 0.440 1.235 ;
        RECT  0.070 1.050 0.210 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.320 -0.210 0.840 0.210 ;
        RECT  0.150 -0.210 0.320 0.890 ;
        RECT  0.000 -0.210 0.150 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.320 2.310 0.840 2.730 ;
        RECT  0.150 1.525 0.320 2.730 ;
        RECT  0.000 2.310 0.150 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 0.840 2.520 ;
	 END
END INVX1AD
MACRO INVX20AD
    CLASS CORE ;
    FOREIGN INVX20AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.355 0.400 3.525 2.120 ;
        RECT  2.805 0.940 3.355 1.690 ;
        RECT  2.635 0.400 2.805 2.120 ;
        RECT  2.085 0.890 2.635 1.690 ;
        RECT  1.915 0.395 2.085 2.150 ;
        RECT  1.685 0.645 1.915 1.690 ;
        RECT  1.390 0.645 1.685 0.900 ;
        RECT  1.390 1.360 1.685 1.690 ;
        RECT  1.170 0.375 1.390 0.900 ;
        RECT  1.170 1.360 1.390 2.165 ;
        RECT  0.670 0.645 1.170 0.900 ;
        RECT  0.670 1.360 1.170 1.690 ;
        RECT  0.450 0.375 0.670 0.900 ;
        RECT  0.460 1.360 0.670 2.145 ;
        END
        AntennaDiffArea 2.11 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.070 1.560 1.190 ;
        RECT  0.070 1.070 0.210 1.445 ;
        END
        AntennaGateArea 1.62 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.930 -0.210 4.200 0.210 ;
        RECT  3.670 -0.210 3.930 0.785 ;
        RECT  3.190 -0.210 3.670 0.210 ;
        RECT  2.970 -0.210 3.190 0.785 ;
        RECT  2.490 -0.210 2.970 0.210 ;
        RECT  2.230 -0.210 2.490 0.760 ;
        RECT  1.770 -0.210 2.230 0.210 ;
        RECT  1.510 -0.210 1.770 0.525 ;
        RECT  1.050 -0.210 1.510 0.210 ;
        RECT  0.790 -0.210 1.050 0.525 ;
        RECT  0.285 -0.210 0.790 0.210 ;
        RECT  0.115 -0.210 0.285 0.785 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.885 2.310 4.200 2.730 ;
        RECT  3.715 1.475 3.885 2.730 ;
        RECT  3.190 2.310 3.715 2.730 ;
        RECT  2.970 1.845 3.190 2.730 ;
        RECT  2.470 2.310 2.970 2.730 ;
        RECT  2.250 1.845 2.470 2.730 ;
        RECT  1.750 2.310 2.250 2.730 ;
        RECT  1.530 1.845 1.750 2.730 ;
        RECT  1.030 2.310 1.530 2.730 ;
        RECT  1.005 2.080 1.030 2.730 ;
        RECT  0.835 1.845 1.005 2.730 ;
        RECT  0.810 2.080 0.835 2.730 ;
        RECT  0.285 2.310 0.810 2.730 ;
        RECT  0.115 1.585 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
	 END
END INVX20AD
MACRO INVX2AD
    CLASS CORE ;
    FOREIGN INVX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.715 0.685 0.770 1.565 ;
        RECT  0.600 0.425 0.715 2.075 ;
        RECT  0.545 0.425 0.600 0.855 ;
        RECT  0.545 1.385 0.600 2.075 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.090 0.480 1.265 ;
        RECT  0.070 1.090 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.355 -0.210 0.840 0.210 ;
        RECT  0.185 -0.210 0.355 0.855 ;
        RECT  0.000 -0.210 0.185 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.355 2.310 0.840 2.730 ;
        RECT  0.185 1.585 0.355 2.730 ;
        RECT  0.000 2.310 0.185 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 0.840 2.520 ;
	 END
END INVX2AD
MACRO INVX3AD
    CLASS CORE ;
    FOREIGN INVX3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.390 0.770 2.020 ;
        RECT  0.475 0.390 0.630 0.870 ;
        RECT  0.475 1.500 0.630 2.020 ;
        END
        AntennaDiffArea 0.318 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.305 1.000 0.510 1.375 ;
        RECT  0.130 1.000 0.305 1.260 ;
        END
        AntennaGateArea 0.244 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 -0.210 1.120 0.210 ;
        RECT  0.890 -0.210 1.050 0.890 ;
        RECT  0.285 -0.210 0.890 0.210 ;
        RECT  0.115 -0.210 0.285 0.870 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 2.310 1.120 2.730 ;
        RECT  0.890 1.500 1.050 2.730 ;
        RECT  0.285 2.310 0.890 2.730 ;
        RECT  0.115 1.500 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
	 END
END INVX3AD
MACRO INVX4AD
    CLASS CORE ;
    FOREIGN INVX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 1.005 0.770 1.515 ;
        RECT  0.740 0.685 0.750 1.515 ;
        RECT  0.670 0.685 0.740 2.155 ;
        RECT  0.620 0.330 0.670 2.155 ;
        RECT  0.450 0.330 0.620 0.850 ;
        RECT  0.450 1.635 0.620 2.155 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.040 0.490 1.300 ;
        RECT  0.110 1.040 0.210 1.655 ;
        RECT  0.070 1.130 0.110 1.655 ;
        END
        AntennaGateArea 0.3249 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.030 -0.210 1.120 0.210 ;
        RECT  0.870 -0.210 1.030 0.850 ;
        RECT  0.280 -0.210 0.870 0.210 ;
        RECT  0.105 -0.210 0.280 0.850 ;
        RECT  0.000 -0.210 0.105 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.025 2.310 1.120 2.730 ;
        RECT  0.860 1.635 1.025 2.730 ;
        RECT  0.290 2.310 0.860 2.730 ;
        RECT  0.110 1.775 0.290 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
	 END
END INVX4AD
MACRO INVX5AD
    CLASS CORE ;
    FOREIGN INVX5AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.370 1.330 2.120 ;
        RECT  0.445 0.645 1.170 0.815 ;
        RECT  0.445 1.555 1.170 1.725 ;
        END
        AntennaDiffArea 0.712 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.270 1.030 0.770 1.375 ;
        END
        AntennaGateArea 0.4044 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 -0.210 1.400 0.210 ;
        RECT  0.670 -0.210 0.930 0.290 ;
        RECT  0.255 -0.210 0.670 0.210 ;
        RECT  0.085 -0.210 0.255 0.815 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.930 2.310 1.400 2.730 ;
        RECT  0.670 2.090 0.930 2.730 ;
        RECT  0.255 2.310 0.670 2.730 ;
        RECT  0.085 1.555 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
	 END
END INVX5AD
MACRO INVX6AD
    CLASS CORE ;
    FOREIGN INVX6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.410 0.395 1.535 0.950 ;
        RECT  1.410 1.550 1.515 1.980 ;
        RECT  1.355 0.395 1.410 1.980 ;
        RECT  1.345 0.770 1.355 1.980 ;
        RECT  1.035 0.770 1.345 1.730 ;
        RECT  0.730 0.770 1.035 0.950 ;
        RECT  0.725 1.550 1.035 1.730 ;
        RECT  0.550 0.395 0.730 0.950 ;
        RECT  0.545 1.550 0.725 1.980 ;
        END
        AntennaDiffArea 0.831 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.070 0.850 1.375 ;
        END
        AntennaGateArea 0.486 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.175 -0.210 1.680 0.210 ;
        RECT  0.915 -0.210 1.175 0.650 ;
        RECT  0.370 -0.210 0.915 0.210 ;
        RECT  0.170 -0.210 0.370 0.875 ;
        RECT  0.000 -0.210 0.170 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.170 2.310 1.680 2.730 ;
        RECT  0.910 1.870 1.170 2.730 ;
        RECT  0.380 2.310 0.910 2.730 ;
        RECT  0.355 1.590 0.380 2.730 ;
        RECT  0.185 1.565 0.355 2.730 ;
        RECT  0.160 1.590 0.185 2.730 ;
        RECT  0.000 2.310 0.160 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
	 END
END INVX6AD
MACRO INVX8AD
    CLASS CORE ;
    FOREIGN INVX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.295 0.475 1.495 2.190 ;
        RECT  1.045 0.795 1.295 1.710 ;
        RECT  0.750 0.795 1.045 0.995 ;
        RECT  0.730 1.460 1.045 1.710 ;
        RECT  0.550 0.475 0.750 0.995 ;
        RECT  0.470 1.460 0.730 2.190 ;
        END
        AntennaDiffArea 0.914 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.120 0.840 1.240 ;
        RECT  0.070 1.120 0.210 1.375 ;
        END
        AntennaGateArea 0.648 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.835 -0.210 1.960 0.210 ;
        RECT  1.665 -0.210 1.835 0.690 ;
        RECT  1.100 -0.210 1.665 0.210 ;
        RECT  0.920 -0.210 1.100 0.675 ;
        RECT  0.375 -0.210 0.920 0.210 ;
        RECT  0.205 -0.210 0.375 0.695 ;
        RECT  0.000 -0.210 0.205 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.835 2.310 1.960 2.730 ;
        RECT  1.665 1.500 1.835 2.730 ;
        RECT  1.125 2.310 1.665 2.730 ;
        RECT  0.865 1.830 1.125 2.730 ;
        RECT  0.295 2.310 0.865 2.730 ;
        RECT  0.125 1.500 0.295 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
	 END
END INVX8AD
MACRO INVXLAD
    CLASS CORE ;
    FOREIGN INVXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 0.735 0.770 1.710 ;
        RECT  0.510 0.735 0.610 0.905 ;
        RECT  0.510 1.540 0.610 1.710 ;
        END
        AntennaDiffArea 0.144 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.070 0.465 1.235 ;
        RECT  0.070 1.070 0.210 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.320 -0.210 0.840 0.210 ;
        RECT  0.150 -0.210 0.320 0.905 ;
        RECT  0.000 -0.210 0.150 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.320 2.310 0.840 2.730 ;
        RECT  0.150 1.495 0.320 2.730 ;
        RECT  0.000 2.310 0.150 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 0.840 2.520 ;
	 END
END INVXLAD
MACRO MDFFHQX1AD
    CLASS CORE ;
    FOREIGN MDFFHQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 0.790 1.610 1.310 ;
        END
        AntennaGateArea 0.098 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.025 1.425 8.050 1.655 ;
        RECT  8.000 0.400 8.025 0.570 ;
        RECT  8.000 1.425 8.025 2.030 ;
        RECT  7.880 0.400 8.000 2.030 ;
        RECT  7.855 0.400 7.880 0.570 ;
        RECT  7.855 1.560 7.880 2.030 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.890 1.195 ;
        END
        AntennaGateArea 0.049 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.220 0.860 2.490 1.135 ;
        END
        AntennaGateArea 0.049 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.870 0.910 3.010 1.375 ;
        END
        AntennaGateArea 0.114 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.640 -0.210 8.120 0.210 ;
        RECT  7.470 -0.210 7.640 0.370 ;
        RECT  7.150 -0.210 7.470 0.210 ;
        RECT  6.980 -0.210 7.150 0.370 ;
        RECT  5.610 -0.210 6.980 0.210 ;
        RECT  5.440 -0.210 5.610 0.280 ;
        RECT  4.355 -0.210 5.440 0.210 ;
        RECT  4.185 -0.210 4.355 0.270 ;
        RECT  3.675 -0.210 4.185 0.210 ;
        RECT  3.505 -0.210 3.675 0.755 ;
        RECT  2.595 -0.210 3.505 0.210 ;
        RECT  2.425 -0.210 2.595 0.325 ;
        RECT  0.985 -0.210 2.425 0.210 ;
        RECT  0.815 -0.210 0.985 0.705 ;
        RECT  0.000 -0.210 0.815 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.665 2.310 8.120 2.730 ;
        RECT  7.495 1.560 7.665 2.730 ;
        RECT  7.010 2.310 7.495 2.730 ;
        RECT  6.840 1.825 7.010 2.730 ;
        RECT  5.610 2.310 6.840 2.730 ;
        RECT  5.440 2.265 5.610 2.730 ;
        RECT  4.425 2.310 5.440 2.730 ;
        RECT  4.255 2.265 4.425 2.730 ;
        RECT  3.105 2.310 4.255 2.730 ;
        RECT  2.935 2.265 3.105 2.730 ;
        RECT  2.465 2.310 2.935 2.730 ;
        RECT  2.295 2.265 2.465 2.730 ;
        RECT  1.045 2.310 2.295 2.730 ;
        RECT  0.875 2.265 1.045 2.730 ;
        RECT  0.000 2.310 0.875 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.120 2.520 ;
        LAYER M1 ;
        RECT  7.720 0.830 7.760 1.350 ;
        RECT  7.600 0.500 7.720 1.350 ;
        RECT  6.875 0.500 7.600 0.620 ;
        RECT  7.360 0.740 7.480 1.000 ;
        RECT  7.285 0.830 7.360 1.000 ;
        RECT  7.115 0.830 7.285 1.645 ;
        RECT  6.840 1.160 7.115 1.330 ;
        RECT  6.755 0.500 6.875 0.710 ;
        RECT  6.350 0.590 6.755 0.710 ;
        RECT  6.655 0.850 6.680 1.090 ;
        RECT  6.535 0.850 6.655 2.190 ;
        RECT  6.510 0.850 6.535 1.090 ;
        RECT  6.485 1.980 6.535 2.190 ;
        RECT  5.195 1.980 6.485 2.100 ;
        RECT  6.230 0.590 6.350 1.750 ;
        RECT  6.090 0.330 6.275 0.450 ;
        RECT  6.180 0.685 6.230 0.855 ;
        RECT  6.180 1.580 6.230 1.750 ;
        RECT  5.970 0.330 6.090 0.540 ;
        RECT  5.915 0.665 6.035 1.750 ;
        RECT  5.220 0.420 5.970 0.540 ;
        RECT  5.775 0.665 5.915 0.905 ;
        RECT  5.820 1.580 5.915 1.750 ;
        RECT  5.660 1.045 5.780 1.360 ;
        RECT  5.530 0.785 5.775 0.905 ;
        RECT  5.015 1.240 5.660 1.360 ;
        RECT  5.360 0.785 5.530 1.120 ;
        RECT  5.270 0.950 5.360 1.120 ;
        RECT  4.960 0.355 5.220 0.540 ;
        RECT  5.145 1.980 5.195 2.185 ;
        RECT  5.025 1.735 5.145 2.185 ;
        RECT  4.965 0.665 5.060 0.785 ;
        RECT  4.720 1.735 5.025 1.855 ;
        RECT  4.965 1.240 5.015 1.615 ;
        RECT  4.845 0.665 4.965 1.615 ;
        RECT  4.140 0.420 4.960 0.540 ;
        RECT  4.620 2.020 4.880 2.180 ;
        RECT  4.800 0.665 4.845 0.785 ;
        RECT  4.600 0.890 4.720 1.855 ;
        RECT  1.850 2.020 4.620 2.140 ;
        RECT  4.280 0.890 4.600 1.010 ;
        RECT  3.790 1.735 4.600 1.855 ;
        RECT  4.360 1.150 4.480 1.410 ;
        RECT  4.140 1.245 4.360 1.365 ;
        RECT  4.060 0.420 4.140 1.365 ;
        RECT  4.020 0.420 4.060 1.560 ;
        RECT  3.865 0.575 4.020 0.745 ;
        RECT  3.800 1.245 4.020 1.560 ;
        RECT  3.315 0.890 3.900 1.010 ;
        RECT  3.615 1.245 3.800 1.365 ;
        RECT  3.530 1.735 3.790 1.900 ;
        RECT  3.445 1.195 3.615 1.365 ;
        RECT  2.330 1.735 3.530 1.855 ;
        RECT  3.195 0.585 3.315 1.615 ;
        RECT  3.145 0.585 3.195 0.755 ;
        RECT  2.630 1.495 3.195 1.615 ;
        RECT  2.750 0.595 2.975 0.765 ;
        RECT  2.630 0.595 2.750 1.375 ;
        RECT  2.330 1.255 2.630 1.375 ;
        RECT  2.210 1.255 2.330 1.855 ;
        RECT  2.090 0.620 2.290 0.740 ;
        RECT  1.970 0.620 2.090 1.725 ;
        RECT  1.730 0.550 1.850 2.140 ;
        RECT  1.585 1.525 1.730 1.695 ;
        RECT  0.205 2.020 1.730 2.140 ;
        RECT  1.565 0.330 1.615 0.500 ;
        RECT  1.445 0.330 1.565 0.590 ;
        RECT  1.345 0.470 1.445 0.590 ;
        RECT  1.295 1.445 1.395 1.615 ;
        RECT  1.295 0.470 1.345 0.705 ;
        RECT  1.175 0.470 1.295 1.860 ;
        RECT  0.590 1.740 1.175 1.860 ;
        RECT  0.505 1.400 0.640 1.570 ;
        RECT  0.505 0.535 0.625 0.705 ;
        RECT  0.330 1.740 0.590 1.890 ;
        RECT  0.385 0.535 0.505 1.570 ;
        RECT  0.205 0.535 0.265 0.705 ;
        RECT  0.205 1.415 0.265 1.585 ;
        RECT  0.085 0.535 0.205 2.140 ;
    END
END MDFFHQX1AD
MACRO MDFFHQX2AD
    CLASS CORE ;
    FOREIGN MDFFHQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.205 0.770 1.375 0.980 ;
        RECT  0.770 0.860 1.205 0.980 ;
        RECT  0.600 0.860 0.770 1.120 ;
        END
        AntennaGateArea 0.125 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.210 0.360 8.330 2.155 ;
        RECT  8.160 0.360 8.210 0.920 ;
        RECT  8.160 1.375 8.210 2.155 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.110 1.350 1.375 ;
        RECT  0.890 1.110 1.190 1.270 ;
        END
        AntennaGateArea 0.077 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.840 2.505 1.140 ;
        END
        AntennaGateArea 0.077 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.870 0.935 3.010 1.375 ;
        END
        AntennaGateArea 0.117 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.795 -0.210 8.400 0.210 ;
        RECT  7.625 -0.210 7.795 0.255 ;
        RECT  5.810 -0.210 7.625 0.210 ;
        RECT  5.640 -0.210 5.810 0.255 ;
        RECT  4.445 -0.210 5.640 0.210 ;
        RECT  4.275 -0.210 4.445 0.255 ;
        RECT  3.315 -0.210 4.275 0.210 ;
        RECT  3.145 -0.210 3.315 0.325 ;
        RECT  2.715 -0.210 3.145 0.210 ;
        RECT  2.545 -0.210 2.715 0.420 ;
        RECT  1.215 -0.210 2.545 0.210 ;
        RECT  1.045 -0.210 1.215 0.630 ;
        RECT  0.000 -0.210 1.045 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.955 2.310 8.400 2.730 ;
        RECT  7.795 1.385 7.955 2.730 ;
        RECT  7.310 2.310 7.795 2.730 ;
        RECT  7.310 1.340 7.435 1.600 ;
        RECT  7.190 1.340 7.310 2.730 ;
        RECT  6.015 2.310 7.190 2.730 ;
        RECT  5.895 2.190 6.015 2.730 ;
        RECT  4.525 2.310 5.895 2.730 ;
        RECT  4.355 2.265 4.525 2.730 ;
        RECT  3.215 2.310 4.355 2.730 ;
        RECT  3.045 2.265 3.215 2.730 ;
        RECT  2.645 2.310 3.045 2.730 ;
        RECT  2.475 2.265 2.645 2.730 ;
        RECT  1.235 2.310 2.475 2.730 ;
        RECT  1.065 2.265 1.235 2.730 ;
        RECT  0.000 2.310 1.065 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.400 2.520 ;
        LAYER M1 ;
        RECT  8.025 1.045 8.075 1.215 ;
        RECT  7.905 0.380 8.025 1.215 ;
        RECT  6.810 0.380 7.905 0.500 ;
        RECT  7.635 1.005 7.675 1.980 ;
        RECT  7.555 0.725 7.635 1.980 ;
        RECT  7.465 0.725 7.555 1.175 ;
        RECT  7.430 1.720 7.555 1.980 ;
        RECT  7.195 1.005 7.465 1.175 ;
        RECT  7.050 0.630 7.190 0.750 ;
        RECT  7.050 1.890 7.070 2.150 ;
        RECT  6.930 0.630 7.050 2.150 ;
        RECT  5.755 1.925 6.930 2.045 ;
        RECT  6.690 0.380 6.810 1.780 ;
        RECT  6.650 0.380 6.690 0.640 ;
        RECT  6.645 1.520 6.690 1.780 ;
        RECT  6.520 0.800 6.570 1.060 ;
        RECT  6.400 0.380 6.520 1.060 ;
        RECT  6.300 1.375 6.470 1.805 ;
        RECT  5.345 0.380 6.400 0.500 ;
        RECT  6.270 1.375 6.300 1.545 ;
        RECT  6.150 0.620 6.270 1.545 ;
        RECT  6.100 0.620 6.150 0.790 ;
        RECT  5.670 0.620 6.100 0.740 ;
        RECT  5.950 0.880 6.020 1.140 ;
        RECT  5.830 0.880 5.950 1.425 ;
        RECT  5.315 1.305 5.830 1.425 ;
        RECT  5.615 1.925 5.755 2.180 ;
        RECT  5.550 0.620 5.670 1.120 ;
        RECT  5.495 1.770 5.615 2.180 ;
        RECT  5.500 0.950 5.550 1.120 ;
        RECT  4.930 1.770 5.495 1.890 ;
        RECT  5.205 2.020 5.375 2.190 ;
        RECT  5.085 0.345 5.345 0.500 ;
        RECT  5.225 1.305 5.315 1.620 ;
        RECT  5.105 0.625 5.225 1.620 ;
        RECT  1.870 2.020 5.205 2.140 ;
        RECT  4.965 0.625 5.105 0.745 ;
        RECT  4.255 0.380 5.085 0.500 ;
        RECT  4.810 0.960 4.930 1.890 ;
        RECT  4.625 0.960 4.810 1.080 ;
        RECT  3.845 1.770 4.810 1.890 ;
        RECT  4.550 1.270 4.670 1.530 ;
        RECT  4.455 0.910 4.625 1.080 ;
        RECT  4.255 1.340 4.550 1.460 ;
        RECT  4.135 0.380 4.255 1.575 ;
        RECT  3.895 0.575 4.135 0.745 ;
        RECT  3.955 1.340 4.135 1.575 ;
        RECT  3.705 0.915 3.995 1.035 ;
        RECT  3.770 1.340 3.955 1.460 ;
        RECT  3.675 1.720 3.845 1.890 ;
        RECT  3.510 1.225 3.770 1.460 ;
        RECT  3.535 0.590 3.705 1.035 ;
        RECT  2.610 1.770 3.675 1.890 ;
        RECT  3.250 0.915 3.535 1.035 ;
        RECT  3.130 0.915 3.250 1.620 ;
        RECT  2.750 1.500 3.130 1.620 ;
        RECT  2.835 0.600 3.005 0.770 ;
        RECT  2.750 0.650 2.835 0.770 ;
        RECT  2.630 0.650 2.750 1.380 ;
        RECT  2.610 1.260 2.630 1.380 ;
        RECT  2.490 1.260 2.610 1.890 ;
        RECT  2.190 0.515 2.325 0.685 ;
        RECT  2.190 1.540 2.255 1.710 ;
        RECT  2.070 0.515 2.190 1.710 ;
        RECT  1.870 0.480 1.940 1.280 ;
        RECT  1.820 0.480 1.870 2.140 ;
        RECT  1.750 1.160 1.820 2.140 ;
        RECT  0.495 2.020 1.750 2.140 ;
        RECT  1.630 0.780 1.690 1.040 ;
        RECT  1.555 0.460 1.630 1.620 ;
        RECT  1.510 0.460 1.555 1.855 ;
        RECT  1.405 0.460 1.510 0.630 ;
        RECT  1.385 1.500 1.510 1.855 ;
        RECT  1.070 1.500 1.385 1.620 ;
        RECT  0.950 1.390 1.070 1.620 ;
        RECT  0.740 1.390 0.950 1.510 ;
        RECT  0.685 0.445 0.855 0.740 ;
        RECT  0.830 1.715 0.855 1.885 ;
        RECT  0.685 1.630 0.830 1.885 ;
        RECT  0.600 1.250 0.740 1.510 ;
        RECT  0.470 0.620 0.685 0.740 ;
        RECT  0.470 1.630 0.685 1.750 ;
        RECT  0.220 0.380 0.540 0.500 ;
        RECT  0.325 1.870 0.495 2.140 ;
        RECT  0.350 0.620 0.470 1.750 ;
        RECT  0.220 1.870 0.325 1.990 ;
        RECT  0.100 0.380 0.220 1.990 ;
    END
END MDFFHQX2AD
MACRO MDFFHQX4AD
    CLASS CORE ;
    FOREIGN MDFFHQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.775 1.160 1.035 ;
        RECT  0.490 0.865 1.040 1.035 ;
        RECT  0.350 0.865 0.490 1.160 ;
        END
        AntennaGateArea 0.191 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.025 1.005 11.130 1.515 ;
        RECT  10.855 0.420 11.025 2.130 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.675 1.165 1.095 1.335 ;
        END
        AntennaGateArea 0.143 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.585 2.730 1.095 ;
        RECT  2.530 0.770 2.590 1.095 ;
        RECT  2.410 0.770 2.530 1.195 ;
        END
        AntennaGateArea 0.143 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.365 1.055 3.535 1.225 ;
        RECT  3.105 0.910 3.365 1.330 ;
        END
        AntennaGateArea 0.191 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.385 -0.210 11.480 0.210 ;
        RECT  11.215 -0.210 11.385 0.810 ;
        RECT  10.665 -0.210 11.215 0.210 ;
        RECT  10.495 -0.210 10.665 0.535 ;
        RECT  10.085 -0.210 10.495 0.210 ;
        RECT  9.915 -0.210 10.085 0.255 ;
        RECT  8.050 -0.210 9.915 0.210 ;
        RECT  7.880 -0.210 8.050 0.255 ;
        RECT  7.195 -0.210 7.880 0.210 ;
        RECT  7.025 -0.210 7.195 0.255 ;
        RECT  5.995 -0.210 7.025 0.210 ;
        RECT  5.825 -0.210 5.995 0.255 ;
        RECT  4.695 -0.210 5.825 0.210 ;
        RECT  4.525 -0.210 4.695 0.360 ;
        RECT  3.415 -0.210 4.525 0.210 ;
        RECT  3.245 -0.210 3.415 0.745 ;
        RECT  2.785 -0.210 3.245 0.210 ;
        RECT  2.615 -0.210 2.785 0.255 ;
        RECT  1.255 -0.210 2.615 0.210 ;
        RECT  0.825 -0.210 1.255 0.255 ;
        RECT  0.000 -0.210 0.825 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.385 2.310 11.480 2.730 ;
        RECT  11.215 1.655 11.385 2.730 ;
        RECT  10.665 2.310 11.215 2.730 ;
        RECT  10.495 1.655 10.665 2.730 ;
        RECT  9.985 2.310 10.495 2.730 ;
        RECT  9.725 1.625 9.985 2.730 ;
        RECT  7.995 2.310 9.725 2.730 ;
        RECT  7.825 2.265 7.995 2.730 ;
        RECT  7.235 2.310 7.825 2.730 ;
        RECT  7.065 2.265 7.235 2.730 ;
        RECT  6.405 2.310 7.065 2.730 ;
        RECT  6.235 2.265 6.405 2.730 ;
        RECT  5.095 2.310 6.235 2.730 ;
        RECT  4.925 2.265 5.095 2.730 ;
        RECT  4.295 2.310 4.925 2.730 ;
        RECT  4.125 2.265 4.295 2.730 ;
        RECT  3.395 2.310 4.125 2.730 ;
        RECT  3.225 2.265 3.395 2.730 ;
        RECT  2.815 2.310 3.225 2.730 ;
        RECT  2.645 2.265 2.815 2.730 ;
        RECT  1.455 2.310 2.645 2.730 ;
        RECT  1.285 2.265 1.455 2.730 ;
        RECT  0.000 2.310 1.285 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.480 2.520 ;
        LAYER M1 ;
        RECT  10.565 0.760 10.685 1.505 ;
        RECT  10.055 0.760 10.565 0.880 ;
        RECT  10.320 1.385 10.565 1.505 ;
        RECT  10.055 1.005 10.435 1.265 ;
        RECT  10.150 1.385 10.320 1.770 ;
        RECT  9.790 1.385 10.150 1.505 ;
        RECT  9.890 1.005 10.055 1.125 ;
        RECT  9.770 0.380 9.890 1.125 ;
        RECT  9.620 1.255 9.790 1.505 ;
        RECT  9.225 0.380 9.770 0.500 ;
        RECT  9.480 0.660 9.590 0.920 ;
        RECT  9.360 0.660 9.480 2.100 ;
        RECT  6.775 1.980 9.360 2.100 ;
        RECT  9.145 0.380 9.225 1.550 ;
        RECT  9.105 0.380 9.145 1.735 ;
        RECT  8.530 0.380 9.105 0.500 ;
        RECT  8.975 1.430 9.105 1.735 ;
        RECT  8.835 0.630 8.975 0.750 ;
        RECT  8.210 1.430 8.975 1.550 ;
        RECT  8.715 0.630 8.835 1.270 ;
        RECT  8.615 1.690 8.785 1.860 ;
        RECT  7.670 1.150 8.715 1.270 ;
        RECT  7.670 1.690 8.615 1.810 ;
        RECT  8.360 0.340 8.530 0.770 ;
        RECT  8.015 0.890 8.355 1.010 ;
        RECT  7.895 0.380 8.015 1.010 ;
        RECT  4.965 0.380 7.895 0.500 ;
        RECT  7.615 0.635 7.670 1.810 ;
        RECT  7.550 0.635 7.615 1.860 ;
        RECT  7.500 0.635 7.550 0.805 ;
        RECT  7.445 1.345 7.550 1.860 ;
        RECT  7.090 1.345 7.445 1.465 ;
        RECT  7.380 0.945 7.420 1.205 ;
        RECT  7.260 0.620 7.380 1.205 ;
        RECT  6.655 0.620 7.260 0.740 ;
        RECT  6.970 0.900 7.090 1.465 ;
        RECT  6.655 1.760 6.775 2.100 ;
        RECT  6.535 0.620 6.655 1.590 ;
        RECT  6.605 1.760 6.655 1.930 ;
        RECT  5.485 1.760 6.605 1.880 ;
        RECT  6.350 0.620 6.535 0.780 ;
        RECT  6.485 1.385 6.535 1.590 ;
        RECT  5.775 1.470 6.485 1.590 ;
        RECT  5.130 0.620 6.350 0.740 ;
        RECT  5.400 2.020 5.920 2.190 ;
        RECT  5.485 0.865 5.900 0.985 ;
        RECT  5.605 1.420 5.775 1.590 ;
        RECT  5.365 0.865 5.485 1.880 ;
        RECT  2.050 2.020 5.400 2.140 ;
        RECT  4.835 0.865 5.365 0.985 ;
        RECT  2.770 1.760 5.365 1.880 ;
        RECT  5.100 1.110 5.240 1.230 ;
        RECT  4.980 1.110 5.100 1.620 ;
        RECT  4.315 1.500 4.980 1.620 ;
        RECT  4.845 0.380 4.965 0.610 ;
        RECT  4.315 0.490 4.845 0.610 ;
        RECT  4.665 0.815 4.835 0.985 ;
        RECT  4.195 0.440 4.315 1.620 ;
        RECT  4.145 0.440 4.195 0.610 ;
        RECT  4.025 1.115 4.195 1.285 ;
        RECT  3.805 0.755 4.055 0.925 ;
        RECT  3.685 0.605 3.805 1.620 ;
        RECT  3.605 0.605 3.685 0.775 ;
        RECT  2.890 1.500 3.685 1.620 ;
        RECT  2.985 0.605 3.055 0.775 ;
        RECT  2.865 0.605 2.985 1.350 ;
        RECT  2.770 1.230 2.865 1.350 ;
        RECT  2.650 1.230 2.770 1.880 ;
        RECT  2.290 1.455 2.435 1.885 ;
        RECT  2.290 0.440 2.370 0.610 ;
        RECT  2.170 0.440 2.290 1.885 ;
        RECT  1.930 0.385 2.050 2.140 ;
        RECT  1.835 0.385 1.930 0.815 ;
        RECT  0.255 2.020 1.930 2.140 ;
        RECT  1.680 0.955 1.800 1.215 ;
        RECT  1.680 1.450 1.710 1.710 ;
        RECT  1.560 0.465 1.680 1.860 ;
        RECT  1.520 0.465 1.560 0.725 ;
        RECT  0.920 1.740 1.560 1.860 ;
        RECT  1.280 0.495 1.400 1.620 ;
        RECT  0.615 0.495 1.280 0.615 ;
        RECT  0.525 1.500 1.280 1.620 ;
        RECT  0.660 1.740 0.920 1.900 ;
        RECT  0.445 0.470 0.615 0.640 ;
        RECT  0.205 1.450 0.255 2.140 ;
        RECT  0.205 0.360 0.230 0.880 ;
        RECT  0.085 0.360 0.205 2.140 ;
    END
END MDFFHQX4AD
MACRO MDFFHQX8AD
    CLASS CORE ;
    FOREIGN MDFFHQX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.865 3.290 1.335 ;
        RECT  2.860 1.165 3.150 1.335 ;
        END
        AntennaGateArea 0.345 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.185 0.400 16.355 2.145 ;
        RECT  15.635 1.005 16.185 1.515 ;
        RECT  15.465 0.400 15.635 2.145 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 0.910 0.535 1.175 ;
        END
        AntennaGateArea 0.274 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.945 0.910 4.455 1.165 ;
        END
        AntennaGateArea 0.274 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.100 0.905 6.695 1.075 ;
        END
        AntennaGateArea 0.344 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.715 -0.210 16.800 0.210 ;
        RECT  16.545 -0.210 16.715 0.795 ;
        RECT  15.995 -0.210 16.545 0.210 ;
        RECT  15.825 -0.210 15.995 0.795 ;
        RECT  15.075 -0.210 15.825 0.210 ;
        RECT  14.905 -0.210 15.075 0.255 ;
        RECT  12.355 -0.210 14.905 0.210 ;
        RECT  12.185 -0.210 12.355 0.255 ;
        RECT  11.595 -0.210 12.185 0.210 ;
        RECT  11.425 -0.210 11.595 0.255 ;
        RECT  10.835 -0.210 11.425 0.210 ;
        RECT  10.665 -0.210 10.835 0.255 ;
        RECT  9.930 -0.210 10.665 0.210 ;
        RECT  9.760 -0.210 9.930 0.255 ;
        RECT  8.645 -0.210 9.760 0.210 ;
        RECT  8.385 -0.210 8.645 0.380 ;
        RECT  7.510 -0.210 8.385 0.210 ;
        RECT  7.340 -0.210 7.510 0.255 ;
        RECT  6.735 -0.210 7.340 0.210 ;
        RECT  6.565 -0.210 6.735 0.255 ;
        RECT  5.975 -0.210 6.565 0.210 ;
        RECT  5.805 -0.210 5.975 0.255 ;
        RECT  5.635 -0.210 5.805 0.210 ;
        RECT  5.465 -0.210 5.635 0.255 ;
        RECT  4.690 -0.210 5.465 0.210 ;
        RECT  4.520 -0.210 4.690 0.760 ;
        RECT  3.970 -0.210 4.520 0.210 ;
        RECT  3.800 -0.210 3.970 0.450 ;
        RECT  0.995 -0.210 3.800 0.210 ;
        RECT  0.825 -0.210 0.995 0.255 ;
        RECT  0.255 -0.210 0.825 0.210 ;
        RECT  0.085 -0.210 0.255 0.750 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  16.715 2.310 16.800 2.730 ;
        RECT  16.545 1.445 16.715 2.730 ;
        RECT  15.995 2.310 16.545 2.730 ;
        RECT  15.825 1.785 15.995 2.730 ;
        RECT  15.275 2.310 15.825 2.730 ;
        RECT  15.105 1.835 15.275 2.730 ;
        RECT  14.700 2.310 15.105 2.730 ;
        RECT  14.530 1.725 14.700 2.730 ;
        RECT  12.355 2.310 14.530 2.730 ;
        RECT  12.185 2.265 12.355 2.730 ;
        RECT  11.595 2.310 12.185 2.730 ;
        RECT  11.425 2.265 11.595 2.730 ;
        RECT  10.835 2.310 11.425 2.730 ;
        RECT  10.665 2.265 10.835 2.730 ;
        RECT  9.880 2.310 10.665 2.730 ;
        RECT  9.710 1.930 9.880 2.730 ;
        RECT  8.645 2.310 9.710 2.730 ;
        RECT  8.385 2.130 8.645 2.730 ;
        RECT  7.745 2.310 8.385 2.730 ;
        RECT  7.485 2.130 7.745 2.730 ;
        RECT  6.390 2.310 7.485 2.730 ;
        RECT  6.220 2.265 6.390 2.730 ;
        RECT  5.360 2.310 6.220 2.730 ;
        RECT  5.190 2.265 5.360 2.730 ;
        RECT  4.600 2.310 5.190 2.730 ;
        RECT  4.430 2.265 4.600 2.730 ;
        RECT  3.840 2.310 4.430 2.730 ;
        RECT  3.670 2.265 3.840 2.730 ;
        RECT  0.975 2.310 3.670 2.730 ;
        RECT  0.805 1.755 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.515 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 16.800 2.520 ;
        LAYER M1 ;
        RECT  15.235 1.050 15.285 1.220 ;
        RECT  15.115 0.380 15.235 1.220 ;
        RECT  14.255 0.380 15.115 0.500 ;
        RECT  14.795 0.735 14.965 1.545 ;
        RECT  14.485 1.115 14.795 1.285 ;
        RECT  14.325 0.630 14.495 0.750 ;
        RECT  14.205 0.630 14.325 2.190 ;
        RECT  14.070 0.330 14.255 0.500 ;
        RECT  14.065 2.020 14.205 2.190 ;
        RECT  13.995 0.330 14.070 1.715 ;
        RECT  10.305 2.020 14.065 2.140 ;
        RECT  13.950 0.380 13.995 1.715 ;
        RECT  12.510 0.380 13.950 0.500 ;
        RECT  13.900 1.485 13.950 1.715 ;
        RECT  12.625 1.485 13.900 1.605 ;
        RECT  13.660 0.620 13.830 0.790 ;
        RECT  13.535 1.730 13.705 1.900 ;
        RECT  13.035 0.620 13.660 0.740 ;
        RECT  12.290 1.780 13.535 1.900 ;
        RECT  12.915 0.620 13.035 1.365 ;
        RECT  12.370 0.620 12.915 0.740 ;
        RECT  12.290 1.245 12.915 1.365 ;
        RECT  12.455 1.485 12.625 1.655 ;
        RECT  12.335 0.935 12.505 1.105 ;
        RECT  12.250 0.425 12.370 0.740 ;
        RECT  12.120 0.935 12.335 1.055 ;
        RECT  12.170 1.245 12.290 1.900 ;
        RECT  11.215 0.425 12.250 0.545 ;
        RECT  11.975 1.780 12.170 1.900 ;
        RECT  12.000 0.735 12.120 1.055 ;
        RECT  10.925 0.735 12.000 0.855 ;
        RECT  11.805 1.470 11.975 1.900 ;
        RECT  10.685 0.975 11.875 1.145 ;
        RECT  11.215 1.780 11.805 1.900 ;
        RECT  11.045 0.375 11.215 0.545 ;
        RECT  11.045 1.470 11.215 1.900 ;
        RECT  10.450 1.780 11.045 1.900 ;
        RECT  10.805 0.380 10.925 0.855 ;
        RECT  10.460 0.380 10.805 0.500 ;
        RECT  10.565 0.750 10.685 1.470 ;
        RECT  10.340 0.750 10.565 0.870 ;
        RECT  9.240 1.350 10.565 1.470 ;
        RECT  10.200 0.355 10.460 0.500 ;
        RECT  10.080 0.645 10.340 0.870 ;
        RECT  10.135 1.640 10.305 2.140 ;
        RECT  8.905 0.380 10.200 0.500 ;
        RECT  7.020 1.640 10.135 1.760 ;
        RECT  9.285 0.750 10.080 0.870 ;
        RECT  9.015 2.070 9.415 2.190 ;
        RECT  9.025 0.630 9.285 0.870 ;
        RECT  9.070 1.350 9.240 1.520 ;
        RECT  7.970 1.350 9.070 1.470 ;
        RECT  8.015 0.750 9.025 0.870 ;
        RECT  8.895 1.890 9.015 2.190 ;
        RECT  8.785 0.380 8.905 0.620 ;
        RECT  8.135 1.890 8.895 2.010 ;
        RECT  8.255 0.500 8.785 0.620 ;
        RECT  8.135 0.380 8.255 0.620 ;
        RECT  5.570 0.380 8.135 0.500 ;
        RECT  7.875 1.890 8.135 2.190 ;
        RECT  7.755 0.630 8.015 0.870 ;
        RECT  7.800 1.350 7.970 1.520 ;
        RECT  7.195 1.890 7.875 2.010 ;
        RECT  7.020 0.990 7.800 1.160 ;
        RECT  7.075 1.890 7.195 2.140 ;
        RECT  7.020 0.620 7.175 0.740 ;
        RECT  3.095 2.020 7.075 2.140 ;
        RECT  6.900 0.620 7.020 1.760 ;
        RECT  6.850 1.330 6.900 1.760 ;
        RECT  5.980 0.620 6.400 0.740 ;
        RECT  5.980 1.370 6.080 1.800 ;
        RECT  5.860 0.620 5.980 1.800 ;
        RECT  5.070 0.995 5.860 1.165 ;
        RECT  5.570 1.410 5.740 1.840 ;
        RECT  5.450 0.380 5.570 0.715 ;
        RECT  4.980 1.410 5.570 1.530 ;
        RECT  5.255 0.595 5.450 0.715 ;
        RECT  4.930 0.595 5.255 0.765 ;
        RECT  4.930 1.410 4.980 1.840 ;
        RECT  4.810 0.595 4.930 1.840 ;
        RECT  4.160 0.470 4.330 0.700 ;
        RECT  4.050 1.415 4.220 1.845 ;
        RECT  3.815 0.580 4.160 0.700 ;
        RECT  3.815 1.725 4.050 1.845 ;
        RECT  3.695 0.580 3.815 1.845 ;
        RECT  2.735 1.725 3.695 1.845 ;
        RECT  3.430 0.335 3.550 1.595 ;
        RECT  3.255 0.335 3.430 0.500 ;
        RECT  3.380 1.425 3.430 1.595 ;
        RECT  2.470 0.620 3.275 0.740 ;
        RECT  1.080 0.380 3.255 0.500 ;
        RECT  2.925 1.970 3.095 2.140 ;
        RECT  2.375 2.020 2.925 2.140 ;
        RECT  2.735 0.860 2.895 0.980 ;
        RECT  2.615 0.860 2.735 1.845 ;
        RECT  2.565 1.675 2.615 1.845 ;
        RECT  2.375 0.620 2.470 0.790 ;
        RECT  2.255 0.620 2.375 2.140 ;
        RECT  2.205 1.710 2.255 2.140 ;
        RECT  1.675 2.020 2.205 2.140 ;
        RECT  2.080 0.620 2.130 0.805 ;
        RECT  1.960 0.620 2.080 1.890 ;
        RECT  1.370 0.620 1.960 0.740 ;
        RECT  1.820 1.510 1.960 1.890 ;
        RECT  1.625 0.860 1.795 0.980 ;
        RECT  1.625 1.485 1.675 2.175 ;
        RECT  1.505 0.860 1.625 2.175 ;
        RECT  1.315 0.620 1.370 1.605 ;
        RECT  1.250 0.620 1.315 2.175 ;
        RECT  1.200 0.620 1.250 0.805 ;
        RECT  1.145 1.485 1.250 2.175 ;
        RECT  0.795 1.485 1.145 1.605 ;
        RECT  1.080 1.175 1.130 1.345 ;
        RECT  0.960 0.380 1.080 1.345 ;
        RECT  0.675 0.620 0.795 1.605 ;
        RECT  0.400 0.620 0.675 0.740 ;
        RECT  0.615 1.485 0.675 1.605 ;
        RECT  0.445 1.485 0.615 2.175 ;
    END
END MDFFHQX8AD
MACRO MX2X1AD
    CLASS CORE ;
    FOREIGN MX2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.550 2.450 1.950 ;
        END
        AntennaDiffArea 0.209 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.705 0.375 2.170 ;
        RECT  0.070 1.705 0.115 1.935 ;
        END
        AntennaGateArea 0.1204 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.720 1.145 ;
        END
        AntennaGateArea 0.0724 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.740 0.865 1.925 1.375 ;
        END
        AntennaGateArea 0.072 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.065 -0.210 2.520 0.210 ;
        RECT  1.895 -0.210 2.065 0.745 ;
        RECT  0.625 -0.210 1.895 0.210 ;
        RECT  0.455 -0.210 0.625 0.690 ;
        RECT  0.000 -0.210 0.455 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.090 2.310 2.520 2.730 ;
        RECT  1.830 2.230 2.090 2.730 ;
        RECT  0.665 2.310 1.830 2.730 ;
        RECT  0.495 2.080 0.665 2.730 ;
        RECT  0.000 2.310 0.495 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.050 1.035 2.170 2.000 ;
        RECT  1.320 1.880 2.050 2.000 ;
        RECT  1.620 0.550 1.705 0.720 ;
        RECT  1.620 1.565 1.705 1.735 ;
        RECT  1.500 0.550 1.620 1.735 ;
        RECT  1.200 0.525 1.320 2.000 ;
        RECT  0.940 1.750 1.060 2.150 ;
        RECT  0.840 0.525 0.960 1.630 ;
        RECT  0.720 1.750 0.940 1.870 ;
        RECT  0.600 1.465 0.720 1.870 ;
        RECT  0.265 1.465 0.600 1.585 ;
        RECT  0.215 0.520 0.265 0.690 ;
        RECT  0.215 1.305 0.265 1.585 ;
        RECT  0.095 0.520 0.215 1.585 ;
    END
END MX2X1AD
MACRO MX2X2AD
    CLASS CORE ;
    FOREIGN MX2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 0.370 3.010 2.160 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 2.020 1.690 2.190 ;
        RECT  0.830 2.020 1.430 2.140 ;
        RECT  0.710 1.535 0.830 2.140 ;
        RECT  0.490 1.535 0.710 1.655 ;
        RECT  0.325 0.975 0.490 1.655 ;
        END
        AntennaGateArea 0.1814 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.885 0.770 1.375 ;
        END
        AntennaGateArea 0.129 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.295 0.865 2.450 1.360 ;
        END
        AntennaGateArea 0.1291 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.635 -0.210 3.080 0.210 ;
        RECT  2.465 -0.210 2.635 0.710 ;
        RECT  0.770 -0.210 2.465 0.210 ;
        RECT  0.550 -0.210 0.770 0.485 ;
        RECT  0.000 -0.210 0.550 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.635 2.310 3.080 2.730 ;
        RECT  2.375 2.000 2.635 2.730 ;
        RECT  0.590 2.310 2.375 2.730 ;
        RECT  0.450 1.775 0.590 2.730 ;
        RECT  0.000 2.310 0.450 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  2.595 1.015 2.715 1.870 ;
        RECT  1.750 1.750 2.595 1.870 ;
        RECT  2.175 0.335 2.225 0.765 ;
        RECT  2.175 1.455 2.205 1.625 ;
        RECT  2.055 0.335 2.175 1.625 ;
        RECT  2.025 1.455 2.055 1.625 ;
        RECT  1.815 0.380 1.935 1.095 ;
        RECT  1.045 0.380 1.815 0.500 ;
        RECT  1.705 0.925 1.815 1.095 ;
        RECT  1.575 1.490 1.750 1.870 ;
        RECT  1.575 0.620 1.695 0.790 ;
        RECT  1.455 0.620 1.575 1.870 ;
        RECT  1.285 0.620 1.335 0.790 ;
        RECT  1.165 0.620 1.285 1.760 ;
        RECT  1.070 1.640 1.165 1.760 ;
        RECT  0.950 1.640 1.070 1.900 ;
        RECT  0.925 0.380 1.045 1.380 ;
        RECT  0.265 0.620 0.925 0.740 ;
        RECT  0.205 0.620 0.265 0.850 ;
        RECT  0.205 1.765 0.265 2.025 ;
        RECT  0.085 0.620 0.205 2.025 ;
    END
END MX2X2AD
MACRO MX2X3AD
    CLASS CORE ;
    FOREIGN MX2X3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.915 0.750 3.010 2.190 ;
        RECT  2.860 0.460 2.915 2.190 ;
        RECT  2.745 0.460 2.860 0.890 ;
        RECT  2.770 1.670 2.860 2.190 ;
        END
        AntennaDiffArea 0.318 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 2.020 1.690 2.190 ;
        RECT  0.830 2.020 1.430 2.140 ;
        RECT  0.710 1.535 0.830 2.140 ;
        RECT  0.490 1.535 0.710 1.655 ;
        RECT  0.325 1.020 0.490 1.655 ;
        END
        AntennaGateArea 0.2162 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.910 0.770 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.410 0.865 2.450 1.095 ;
        RECT  2.290 0.865 2.410 1.360 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.250 -0.210 3.360 0.210 ;
        RECT  3.130 -0.210 3.250 0.920 ;
        RECT  2.550 -0.210 3.130 0.210 ;
        RECT  2.390 -0.210 2.550 0.745 ;
        RECT  0.635 -0.210 2.390 0.210 ;
        RECT  0.465 -0.210 0.635 0.525 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.290 2.310 3.360 2.730 ;
        RECT  3.130 1.670 3.290 2.730 ;
        RECT  2.600 2.310 3.130 2.730 ;
        RECT  2.340 2.010 2.600 2.730 ;
        RECT  0.590 2.310 2.340 2.730 ;
        RECT  0.450 1.775 0.590 2.730 ;
        RECT  0.000 2.310 0.450 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.650 1.010 2.740 1.530 ;
        RECT  2.620 1.010 2.650 1.880 ;
        RECT  2.530 1.220 2.620 1.880 ;
        RECT  1.770 1.760 2.530 1.880 ;
        RECT  2.170 1.500 2.240 1.620 ;
        RECT  2.050 0.365 2.170 1.620 ;
        RECT  1.980 1.500 2.050 1.620 ;
        RECT  1.810 0.380 1.930 1.120 ;
        RECT  1.010 0.380 1.810 0.500 ;
        RECT  1.670 1.000 1.810 1.120 ;
        RECT  1.550 1.500 1.770 1.880 ;
        RECT  1.570 0.620 1.690 0.880 ;
        RECT  1.550 0.740 1.570 0.880 ;
        RECT  1.430 0.740 1.550 1.880 ;
        RECT  1.190 0.620 1.310 1.760 ;
        RECT  1.070 1.640 1.190 1.760 ;
        RECT  1.010 1.020 1.070 1.280 ;
        RECT  0.950 1.640 1.070 1.900 ;
        RECT  0.890 0.380 1.010 1.280 ;
        RECT  0.265 0.645 0.890 0.765 ;
        RECT  0.205 0.645 0.265 0.885 ;
        RECT  0.205 1.765 0.265 2.025 ;
        RECT  0.085 0.645 0.205 2.025 ;
    END
END MX2X3AD
MACRO MX2X4AD
    CLASS CORE ;
    FOREIGN MX2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.915 0.655 3.010 2.065 ;
        RECT  2.860 0.390 2.915 2.065 ;
        RECT  2.745 0.390 2.860 0.820 ;
        RECT  2.770 1.545 2.860 2.065 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.430 2.020 1.690 2.190 ;
        RECT  0.830 2.020 1.430 2.140 ;
        RECT  0.710 1.535 0.830 2.140 ;
        RECT  0.490 1.535 0.710 1.655 ;
        RECT  0.325 1.020 0.490 1.655 ;
        END
        AntennaGateArea 0.2162 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.910 0.770 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.410 0.865 2.450 1.095 ;
        RECT  2.290 0.865 2.410 1.360 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.250 -0.210 3.360 0.210 ;
        RECT  3.130 -0.210 3.250 0.850 ;
        RECT  2.555 -0.210 3.130 0.210 ;
        RECT  2.385 -0.210 2.555 0.730 ;
        RECT  0.635 -0.210 2.385 0.210 ;
        RECT  0.465 -0.210 0.635 0.525 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.290 2.310 3.360 2.730 ;
        RECT  3.130 1.495 3.290 2.730 ;
        RECT  2.600 2.310 3.130 2.730 ;
        RECT  2.340 2.010 2.600 2.730 ;
        RECT  0.590 2.310 2.340 2.730 ;
        RECT  0.450 1.775 0.590 2.730 ;
        RECT  0.000 2.310 0.450 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.650 1.025 2.740 1.375 ;
        RECT  2.620 1.025 2.650 1.880 ;
        RECT  2.530 1.190 2.620 1.880 ;
        RECT  1.770 1.760 2.530 1.880 ;
        RECT  2.170 1.500 2.240 1.620 ;
        RECT  2.050 0.365 2.170 1.620 ;
        RECT  1.980 1.500 2.050 1.620 ;
        RECT  1.810 0.380 1.930 1.120 ;
        RECT  1.010 0.380 1.810 0.500 ;
        RECT  1.670 1.000 1.810 1.120 ;
        RECT  1.550 1.500 1.770 1.880 ;
        RECT  1.570 0.620 1.690 0.880 ;
        RECT  1.550 0.740 1.570 0.880 ;
        RECT  1.430 0.740 1.550 1.880 ;
        RECT  1.190 0.620 1.310 1.660 ;
        RECT  1.070 1.540 1.190 1.660 ;
        RECT  1.010 1.020 1.070 1.280 ;
        RECT  0.950 1.540 1.070 1.800 ;
        RECT  0.890 0.380 1.010 1.280 ;
        RECT  0.265 0.645 0.890 0.765 ;
        RECT  0.205 0.645 0.265 0.885 ;
        RECT  0.205 1.765 0.265 2.025 ;
        RECT  0.085 0.645 0.205 2.025 ;
    END
END MX2X4AD
MACRO MX2X6AD
    CLASS CORE ;
    FOREIGN MX2X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.785 3.850 1.690 ;
        RECT  3.700 0.425 3.815 2.150 ;
        RECT  3.645 0.425 3.700 0.925 ;
        RECT  3.645 1.460 3.700 2.150 ;
        RECT  3.095 0.785 3.645 0.925 ;
        RECT  3.095 1.570 3.645 1.750 ;
        RECT  2.925 0.425 3.095 0.925 ;
        RECT  2.925 1.570 3.095 2.075 ;
        END
        AntennaDiffArea 0.795 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 2.020 2.220 2.140 ;
        RECT  0.710 1.535 0.830 2.140 ;
        RECT  0.490 1.535 0.710 1.655 ;
        RECT  0.325 1.020 0.490 1.655 ;
        END
        AntennaGateArea 0.2254 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.910 0.770 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.365 0.865 2.730 1.195 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.500 -0.210 3.920 0.210 ;
        RECT  3.240 -0.210 3.500 0.650 ;
        RECT  2.710 -0.210 3.240 0.210 ;
        RECT  2.540 -0.210 2.710 0.685 ;
        RECT  0.635 -0.210 2.540 0.210 ;
        RECT  0.465 -0.210 0.635 0.525 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.500 2.310 3.920 2.730 ;
        RECT  3.240 1.870 3.500 2.730 ;
        RECT  2.780 2.310 3.240 2.730 ;
        RECT  2.520 2.010 2.780 2.730 ;
        RECT  0.590 2.310 2.520 2.730 ;
        RECT  0.450 1.775 0.590 2.730 ;
        RECT  0.000 2.310 0.450 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  2.970 1.070 3.540 1.240 ;
        RECT  2.850 1.070 2.970 1.450 ;
        RECT  2.710 1.315 2.850 1.450 ;
        RECT  2.590 1.315 2.710 1.880 ;
        RECT  1.550 1.760 2.590 1.880 ;
        RECT  2.245 1.500 2.325 1.620 ;
        RECT  2.125 0.365 2.245 1.620 ;
        RECT  1.805 1.500 2.125 1.620 ;
        RECT  1.885 0.380 2.005 1.280 ;
        RECT  1.010 0.380 1.885 0.500 ;
        RECT  1.550 0.665 1.765 0.835 ;
        RECT  1.430 0.665 1.550 1.880 ;
        RECT  1.190 0.620 1.310 1.760 ;
        RECT  1.070 1.640 1.190 1.760 ;
        RECT  1.010 1.020 1.070 1.280 ;
        RECT  0.950 1.640 1.070 1.900 ;
        RECT  0.890 0.380 1.010 1.280 ;
        RECT  0.265 0.645 0.890 0.765 ;
        RECT  0.205 0.645 0.265 0.885 ;
        RECT  0.205 1.765 0.265 2.025 ;
        RECT  0.085 0.645 0.205 2.025 ;
    END
END MX2X6AD
MACRO MX2X8AD
    CLASS CORE ;
    FOREIGN MX2X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.755 1.000 3.990 1.520 ;
        RECT  3.585 0.385 3.755 2.150 ;
        RECT  3.570 0.785 3.585 1.750 ;
        RECT  3.035 0.785 3.570 0.950 ;
        RECT  3.035 1.570 3.570 1.750 ;
        RECT  2.865 0.390 3.035 0.950 ;
        RECT  2.865 1.570 3.035 2.075 ;
        END
        AntennaDiffArea 0.844 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 2.020 2.220 2.140 ;
        RECT  0.710 1.535 0.830 2.140 ;
        RECT  0.490 1.535 0.710 1.655 ;
        RECT  0.325 1.020 0.490 1.655 ;
        END
        AntennaGateArea 0.2254 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.910 0.770 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.365 0.865 2.730 1.195 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.115 -0.210 4.200 0.210 ;
        RECT  3.945 -0.210 4.115 0.745 ;
        RECT  3.440 -0.210 3.945 0.210 ;
        RECT  3.180 -0.210 3.440 0.650 ;
        RECT  2.650 -0.210 3.180 0.210 ;
        RECT  2.480 -0.210 2.650 0.685 ;
        RECT  0.635 -0.210 2.480 0.210 ;
        RECT  0.465 -0.210 0.635 0.525 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.115 2.310 4.200 2.730 ;
        RECT  3.945 1.845 4.115 2.730 ;
        RECT  3.440 2.310 3.945 2.730 ;
        RECT  3.180 1.870 3.440 2.730 ;
        RECT  2.720 2.310 3.180 2.730 ;
        RECT  2.460 2.010 2.720 2.730 ;
        RECT  0.590 2.310 2.460 2.730 ;
        RECT  0.450 1.775 0.590 2.730 ;
        RECT  0.000 2.310 0.450 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  2.970 1.070 3.280 1.240 ;
        RECT  2.850 1.070 2.970 1.450 ;
        RECT  2.710 1.315 2.850 1.450 ;
        RECT  2.590 1.315 2.710 1.880 ;
        RECT  1.550 1.760 2.590 1.880 ;
        RECT  2.245 1.500 2.325 1.620 ;
        RECT  2.125 0.365 2.245 1.620 ;
        RECT  1.805 1.500 2.125 1.620 ;
        RECT  1.885 0.380 2.005 1.280 ;
        RECT  1.010 0.380 1.885 0.500 ;
        RECT  1.550 0.665 1.765 0.835 ;
        RECT  1.430 0.665 1.550 1.880 ;
        RECT  1.190 0.620 1.310 1.760 ;
        RECT  1.070 1.640 1.190 1.760 ;
        RECT  1.010 1.020 1.070 1.280 ;
        RECT  0.950 1.640 1.070 1.900 ;
        RECT  0.890 0.380 1.010 1.280 ;
        RECT  0.265 0.645 0.890 0.765 ;
        RECT  0.205 0.645 0.265 0.885 ;
        RECT  0.205 1.765 0.265 2.025 ;
        RECT  0.085 0.645 0.205 2.025 ;
    END
END MX2X8AD
MACRO MX2XLAD
    CLASS CORE ;
    FOREIGN MX2XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.460 2.450 1.715 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.705 0.375 2.170 ;
        RECT  0.070 1.705 0.115 1.935 ;
        END
        AntennaGateArea 0.0964 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 0.790 0.720 1.310 ;
        RECT  0.350 0.865 0.600 1.095 ;
        END
        AntennaGateArea 0.0484 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.740 0.865 1.925 1.375 ;
        END
        AntennaGateArea 0.0484 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.110 -0.210 2.520 0.210 ;
        RECT  1.850 -0.210 2.110 0.650 ;
        RECT  0.670 -0.210 1.850 0.210 ;
        RECT  0.410 -0.210 0.670 0.650 ;
        RECT  0.000 -0.210 0.410 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.090 2.310 2.520 2.730 ;
        RECT  1.830 2.120 2.090 2.730 ;
        RECT  0.665 2.310 1.830 2.730 ;
        RECT  0.495 1.990 0.665 2.730 ;
        RECT  0.000 2.310 0.495 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.050 0.790 2.170 2.000 ;
        RECT  1.350 1.880 2.050 2.000 ;
        RECT  1.610 1.510 1.750 1.630 ;
        RECT  1.610 0.505 1.705 0.675 ;
        RECT  1.490 0.505 1.610 1.630 ;
        RECT  1.230 0.505 1.350 2.000 ;
        RECT  1.175 0.505 1.230 0.675 ;
        RECT  1.200 1.360 1.230 1.620 ;
        RECT  0.990 1.750 1.110 2.010 ;
        RECT  0.720 1.750 0.990 1.870 ;
        RECT  0.840 0.460 0.960 1.630 ;
        RECT  0.600 1.465 0.720 1.870 ;
        RECT  0.265 1.465 0.600 1.585 ;
        RECT  0.215 0.505 0.265 0.675 ;
        RECT  0.215 1.415 0.265 1.585 ;
        RECT  0.095 0.505 0.215 1.585 ;
    END
END MX2XLAD
MACRO MX3X1AD
    CLASS CORE ;
    FOREIGN MX3X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.955 0.335 4.970 1.645 ;
        RECT  4.830 0.335 4.955 1.955 ;
        RECT  4.785 0.335 4.830 0.505 ;
        RECT  4.785 1.525 4.830 1.955 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 0.765 3.010 1.285 ;
        END
        AntennaGateArea 0.1414 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 1.890 0.980 2.170 ;
        END
        AntennaGateArea 0.1553 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.170 1.020 0.290 1.375 ;
        RECT  0.070 1.145 0.170 1.375 ;
        END
        AntennaGateArea 0.0724 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.045 1.385 1.215 ;
        RECT  1.160 0.865 1.360 1.215 ;
        END
        AntennaGateArea 0.1044 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.935 2.730 1.375 ;
        END
        AntennaGateArea 0.1074 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.640 -0.210 5.040 0.210 ;
        RECT  4.380 -0.210 4.640 0.390 ;
        RECT  2.825 -0.210 4.380 0.210 ;
        RECT  2.655 -0.210 2.825 0.615 ;
        RECT  1.265 -0.210 2.655 0.210 ;
        RECT  1.095 -0.210 1.265 0.690 ;
        RECT  0.230 -0.210 1.095 0.210 ;
        RECT  0.110 -0.210 0.230 0.420 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.595 2.310 5.040 2.730 ;
        RECT  4.425 1.480 4.595 2.730 ;
        RECT  3.010 2.310 4.425 2.730 ;
        RECT  2.750 2.230 3.010 2.730 ;
        RECT  1.220 2.310 2.750 2.730 ;
        RECT  1.100 1.890 1.220 2.730 ;
        RECT  0.255 2.310 1.100 2.730 ;
        RECT  0.095 1.990 0.255 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.040 2.520 ;
        LAYER M1 ;
        RECT  4.635 0.735 4.705 1.255 ;
        RECT  4.515 0.510 4.635 1.255 ;
        RECT  3.990 0.510 4.515 0.630 ;
        RECT  4.230 0.750 4.395 0.920 ;
        RECT  4.110 0.750 4.230 2.110 ;
        RECT  1.460 1.990 4.110 2.110 ;
        RECT  3.870 0.510 3.990 1.845 ;
        RECT  3.750 1.585 3.870 1.845 ;
        RECT  3.630 0.400 3.750 1.260 ;
        RECT  3.265 0.400 3.630 0.520 ;
        RECT  3.510 1.750 3.580 1.870 ;
        RECT  3.390 0.675 3.510 1.870 ;
        RECT  2.200 1.750 3.390 1.870 ;
        RECT  3.145 0.400 3.265 1.580 ;
        RECT  3.015 0.400 3.145 0.570 ;
        RECT  3.085 1.410 3.145 1.580 ;
        RECT  2.440 1.500 2.650 1.620 ;
        RECT  2.320 0.475 2.440 1.620 ;
        RECT  2.080 0.595 2.200 1.870 ;
        RECT  1.770 0.595 2.080 0.715 ;
        RECT  1.840 0.835 1.960 1.720 ;
        RECT  1.600 0.835 1.840 0.955 ;
        RECT  1.700 1.600 1.840 1.720 ;
        RECT  1.600 1.075 1.720 1.455 ;
        RECT  1.580 1.600 1.700 1.860 ;
        RECT  1.480 0.595 1.600 0.955 ;
        RECT  0.950 1.335 1.600 1.455 ;
        RECT  1.340 1.645 1.460 2.110 ;
        RECT  0.530 1.645 1.340 1.765 ;
        RECT  0.880 1.335 0.950 1.525 ;
        RECT  0.760 0.475 0.880 1.525 ;
        RECT  0.690 1.405 0.760 1.525 ;
        RECT  0.410 0.600 0.530 1.765 ;
    END
END MX3X1AD
MACRO MX3X2AD
    CLASS CORE ;
    FOREIGN MX3X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.490 0.865 5.530 1.095 ;
        RECT  5.370 0.370 5.490 2.180 ;
        RECT  5.330 1.620 5.370 2.180 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.615 1.570 4.970 1.690 ;
        RECT  4.495 1.570 4.615 1.890 ;
        RECT  4.225 1.750 4.495 1.890 ;
        RECT  3.610 1.750 4.225 1.870 ;
        END
        AntennaGateArea 0.2004 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.145 2.730 1.375 ;
        RECT  2.510 1.145 2.630 1.870 ;
        RECT  0.690 1.750 2.510 1.870 ;
        RECT  1.690 0.360 1.950 0.540 ;
        RECT  0.690 0.420 1.690 0.540 ;
        RECT  0.690 1.020 0.805 1.280 ;
        RECT  0.570 0.420 0.690 1.870 ;
        END
        AntennaGateArea 0.2194 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.940 0.210 1.390 ;
        END
        AntennaGateArea 0.13 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.140 1.605 1.375 ;
        END
        AntennaGateArea 0.1619 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 1.010 3.050 1.375 ;
        END
        AntennaGateArea 0.161 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.200 -0.210 5.600 0.210 ;
        RECT  4.940 -0.210 5.200 0.390 ;
        RECT  3.270 -0.210 4.940 0.210 ;
        RECT  3.010 -0.210 3.270 0.390 ;
        RECT  1.295 -0.210 3.010 0.210 ;
        RECT  1.035 -0.210 1.295 0.300 ;
        RECT  0.690 -0.210 1.035 0.210 ;
        RECT  0.430 -0.210 0.690 0.300 ;
        RECT  0.000 -0.210 0.430 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.130 2.310 5.600 2.730 ;
        RECT  5.010 2.060 5.130 2.730 ;
        RECT  3.440 2.310 5.010 2.730 ;
        RECT  3.180 2.230 3.440 2.730 ;
        RECT  1.370 2.310 3.180 2.730 ;
        RECT  1.110 2.230 1.370 2.730 ;
        RECT  0.690 2.310 1.110 2.730 ;
        RECT  0.430 2.230 0.690 2.730 ;
        RECT  0.000 2.310 0.430 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  5.130 0.510 5.250 1.210 ;
        RECT  5.090 1.330 5.210 1.940 ;
        RECT  4.415 0.510 5.130 0.630 ;
        RECT  5.035 1.040 5.130 1.210 ;
        RECT  4.915 1.330 5.090 1.450 ;
        RECT  4.890 1.820 5.090 1.940 ;
        RECT  4.795 0.750 4.915 1.450 ;
        RECT  4.770 1.820 4.890 2.130 ;
        RECT  4.640 0.750 4.795 0.870 ;
        RECT  3.680 2.010 4.770 2.130 ;
        RECT  4.375 0.435 4.415 1.025 ;
        RECT  4.245 0.435 4.375 1.630 ;
        RECT  4.205 1.460 4.245 1.630 ;
        RECT  3.950 0.720 4.060 1.560 ;
        RECT  3.940 0.335 3.950 1.560 ;
        RECT  3.830 0.335 3.940 0.855 ;
        RECT  3.800 1.440 3.940 1.560 ;
        RECT  2.480 0.510 3.830 0.630 ;
        RECT  3.680 0.975 3.820 1.240 ;
        RECT  3.650 0.750 3.680 1.240 ;
        RECT  3.560 1.990 3.680 2.130 ;
        RECT  3.530 0.750 3.650 1.590 ;
        RECT  0.450 1.990 3.560 2.110 ;
        RECT  3.420 0.750 3.530 0.870 ;
        RECT  3.490 1.330 3.530 1.590 ;
        RECT  3.175 0.750 3.295 1.720 ;
        RECT  2.650 0.750 3.175 0.870 ;
        RECT  2.940 1.600 3.175 1.720 ;
        RECT  2.820 1.600 2.940 1.860 ;
        RECT  2.390 0.510 2.480 0.780 ;
        RECT  2.270 0.510 2.390 1.620 ;
        RECT  2.030 0.660 2.150 1.620 ;
        RECT  1.520 0.660 2.030 0.780 ;
        RECT  1.540 1.500 2.030 1.620 ;
        RECT  1.790 0.900 1.910 1.330 ;
        RECT  1.070 0.900 1.790 1.020 ;
        RECT  0.950 0.695 1.070 1.585 ;
        RECT  0.810 0.695 0.950 0.865 ;
        RECT  0.810 1.465 0.950 1.585 ;
        RECT  0.330 0.660 0.450 2.110 ;
        RECT  0.255 0.660 0.330 0.820 ;
        RECT  0.110 1.510 0.330 2.110 ;
        RECT  0.085 0.390 0.255 0.820 ;
    END
END MX3X2AD
MACRO MX3X4AD
    CLASS CORE ;
    FOREIGN MX3X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.705 0.370 5.810 1.655 ;
        RECT  5.670 0.370 5.705 2.160 ;
        RECT  5.560 0.370 5.670 0.890 ;
        RECT  5.535 1.470 5.670 2.160 ;
        END
        AntennaDiffArea 0.438 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.690 1.030 4.800 1.655 ;
        RECT  4.680 1.030 4.690 1.870 ;
        RECT  4.550 1.420 4.680 1.870 ;
        RECT  3.610 1.750 4.550 1.870 ;
        END
        AntennaGateArea 0.2214 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.145 2.730 1.375 ;
        RECT  2.510 1.145 2.630 1.870 ;
        RECT  0.690 1.750 2.510 1.870 ;
        RECT  1.690 0.360 1.950 0.540 ;
        RECT  0.690 0.420 1.690 0.540 ;
        RECT  0.690 1.020 0.805 1.280 ;
        RECT  0.570 0.420 0.690 1.870 ;
        END
        AntennaGateArea 0.2194 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.940 0.210 1.390 ;
        END
        AntennaGateArea 0.162 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.140 1.605 1.375 ;
        END
        AntennaGateArea 0.1619 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 1.010 3.050 1.375 ;
        END
        AntennaGateArea 0.161 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.050 -0.210 6.160 0.210 ;
        RECT  5.930 -0.210 6.050 0.890 ;
        RECT  5.390 -0.210 5.930 0.210 ;
        RECT  5.130 -0.210 5.390 0.390 ;
        RECT  3.270 -0.210 5.130 0.210 ;
        RECT  3.010 -0.210 3.270 0.390 ;
        RECT  1.295 -0.210 3.010 0.210 ;
        RECT  1.035 -0.210 1.295 0.300 ;
        RECT  0.730 -0.210 1.035 0.210 ;
        RECT  0.470 -0.210 0.730 0.300 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.050 2.310 6.160 2.730 ;
        RECT  5.930 1.420 6.050 2.730 ;
        RECT  5.320 2.310 5.930 2.730 ;
        RECT  5.200 1.500 5.320 2.730 ;
        RECT  3.440 2.310 5.200 2.730 ;
        RECT  3.180 2.230 3.440 2.730 ;
        RECT  1.370 2.310 3.180 2.730 ;
        RECT  1.110 2.230 1.370 2.730 ;
        RECT  0.730 2.310 1.110 2.730 ;
        RECT  0.470 2.230 0.730 2.730 ;
        RECT  0.000 2.310 0.470 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.395 1.045 5.445 1.215 ;
        RECT  5.275 0.510 5.395 1.215 ;
        RECT  4.575 0.510 5.275 0.630 ;
        RECT  4.920 0.750 5.040 2.110 ;
        RECT  4.760 0.750 4.920 0.870 ;
        RECT  0.450 1.990 4.920 2.110 ;
        RECT  4.405 0.395 4.575 0.825 ;
        RECT  4.375 0.635 4.405 0.825 ;
        RECT  4.205 0.635 4.375 1.630 ;
        RECT  3.965 0.335 4.085 1.560 ;
        RECT  2.480 0.510 3.965 0.630 ;
        RECT  3.800 1.440 3.965 1.560 ;
        RECT  3.680 0.975 3.845 1.240 ;
        RECT  3.610 0.750 3.680 1.240 ;
        RECT  3.490 0.750 3.610 1.590 ;
        RECT  3.420 0.750 3.490 0.870 ;
        RECT  3.175 0.750 3.295 1.720 ;
        RECT  2.650 0.750 3.175 0.870 ;
        RECT  2.940 1.600 3.175 1.720 ;
        RECT  2.820 1.600 2.940 1.860 ;
        RECT  2.390 0.510 2.480 0.780 ;
        RECT  2.270 0.510 2.390 1.620 ;
        RECT  2.030 0.660 2.150 1.620 ;
        RECT  1.520 0.660 2.030 0.780 ;
        RECT  1.540 1.500 2.030 1.620 ;
        RECT  1.790 0.900 1.910 1.330 ;
        RECT  1.070 0.900 1.790 1.020 ;
        RECT  0.950 0.695 1.070 1.585 ;
        RECT  0.810 0.695 0.950 0.865 ;
        RECT  0.810 1.465 0.950 1.585 ;
        RECT  0.330 0.660 0.450 2.110 ;
        RECT  0.255 0.660 0.330 0.820 ;
        RECT  0.110 1.510 0.330 2.110 ;
        RECT  0.085 0.390 0.255 0.820 ;
    END
END MX3X4AD
MACRO MX3XLAD
    CLASS CORE ;
    FOREIGN MX3XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.830 0.330 4.970 1.825 ;
        RECT  4.785 0.330 4.830 0.500 ;
        RECT  4.785 1.655 4.830 1.825 ;
        END
        AntennaDiffArea 0.143 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 0.780 3.010 1.300 ;
        END
        AntennaGateArea 0.1124 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 1.905 0.980 2.170 ;
        END
        AntennaGateArea 0.1203 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.170 1.020 0.290 1.375 ;
        RECT  0.070 1.145 0.170 1.375 ;
        END
        AntennaGateArea 0.0504 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.045 1.385 1.215 ;
        RECT  1.160 0.865 1.360 1.215 ;
        END
        AntennaGateArea 0.0724 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.935 2.730 1.375 ;
        END
        AntennaGateArea 0.0724 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.620 -0.210 5.040 0.210 ;
        RECT  4.360 -0.210 4.620 0.425 ;
        RECT  2.825 -0.210 4.360 0.210 ;
        RECT  2.655 -0.210 2.825 0.655 ;
        RECT  1.310 -0.210 2.655 0.210 ;
        RECT  1.050 -0.210 1.310 0.730 ;
        RECT  0.230 -0.210 1.050 0.210 ;
        RECT  0.110 -0.210 0.230 0.420 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.595 2.310 5.040 2.730 ;
        RECT  4.425 1.645 4.595 2.730 ;
        RECT  3.010 2.310 4.425 2.730 ;
        RECT  2.750 2.230 3.010 2.730 ;
        RECT  1.220 2.310 2.750 2.730 ;
        RECT  1.100 1.910 1.220 2.730 ;
        RECT  0.255 2.310 1.100 2.730 ;
        RECT  0.095 1.990 0.255 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.040 2.520 ;
        LAYER M1 ;
        RECT  4.660 0.735 4.705 1.255 ;
        RECT  4.540 0.545 4.660 1.255 ;
        RECT  3.990 0.545 4.540 0.665 ;
        RECT  4.230 0.785 4.420 0.905 ;
        RECT  4.110 0.785 4.230 2.110 ;
        RECT  1.460 1.990 4.110 2.110 ;
        RECT  3.870 0.545 3.990 1.860 ;
        RECT  3.725 1.690 3.870 1.860 ;
        RECT  3.630 0.380 3.750 1.385 ;
        RECT  3.255 0.380 3.630 0.500 ;
        RECT  3.510 1.750 3.580 1.870 ;
        RECT  3.390 0.675 3.510 1.870 ;
        RECT  2.200 1.750 3.390 1.870 ;
        RECT  3.135 0.380 3.255 1.570 ;
        RECT  3.015 0.380 3.135 0.655 ;
        RECT  3.085 1.400 3.135 1.570 ;
        RECT  2.440 1.495 2.650 1.615 ;
        RECT  2.320 0.475 2.440 1.615 ;
        RECT  2.080 0.595 2.200 1.870 ;
        RECT  1.770 0.595 2.080 0.715 ;
        RECT  1.840 0.835 1.960 1.695 ;
        RECT  1.600 0.835 1.840 0.955 ;
        RECT  1.700 1.575 1.840 1.695 ;
        RECT  1.600 1.075 1.720 1.455 ;
        RECT  1.580 1.575 1.700 1.860 ;
        RECT  1.480 0.500 1.600 0.955 ;
        RECT  0.950 1.335 1.600 1.455 ;
        RECT  1.340 1.665 1.460 2.110 ;
        RECT  0.530 1.665 1.340 1.785 ;
        RECT  0.880 1.335 0.950 1.545 ;
        RECT  0.760 0.540 0.880 1.545 ;
        RECT  0.690 1.425 0.760 1.545 ;
        RECT  0.410 0.690 0.530 1.785 ;
    END
END MX3XLAD
MACRO MX4X1AD
    CLASS CORE ;
    FOREIGN MX4X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.905 0.595 6.930 1.575 ;
        RECT  6.790 0.595 6.905 1.850 ;
        RECT  6.735 0.595 6.790 0.765 ;
        RECT  6.735 1.420 6.790 1.850 ;
        END
        AntennaDiffArea 0.193 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.200 1.705 6.370 1.935 ;
        RECT  6.080 0.915 6.200 2.140 ;
        RECT  5.430 2.020 6.080 2.140 ;
        RECT  4.910 2.020 5.430 2.190 ;
        END
        AntennaGateArea 0.1494 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.775 1.980 4.035 2.160 ;
        RECT  0.925 1.980 3.775 2.100 ;
        RECT  2.985 0.330 3.285 0.450 ;
        RECT  2.865 0.330 2.985 0.530 ;
        RECT  2.655 0.410 2.865 0.530 ;
        RECT  2.535 0.410 2.655 1.200 ;
        RECT  1.725 0.410 2.535 0.530 ;
        RECT  2.370 1.080 2.535 1.200 ;
        RECT  2.250 1.080 2.370 1.340 ;
        RECT  1.605 0.380 1.725 0.530 ;
        RECT  1.300 0.380 1.605 0.500 ;
        RECT  1.040 0.330 1.300 0.500 ;
        RECT  0.845 0.380 1.040 0.500 ;
        RECT  0.845 1.980 0.925 2.190 ;
        RECT  0.725 0.380 0.845 2.190 ;
        RECT  0.585 2.030 0.725 2.190 ;
        END
        AntennaGateArea 0.2685 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.655 1.890 1.095 ;
        RECT  1.570 0.890 1.750 1.010 ;
        END
        AntennaGateArea 0.1014 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.100 0.865 0.330 1.250 ;
        RECT  0.070 0.865 0.100 1.095 ;
        END
        AntennaGateArea 0.107 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.775 0.910 3.055 1.140 ;
        END
        AntennaGateArea 0.0974 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.270 0.865 4.410 1.230 ;
        RECT  4.205 0.960 4.270 1.230 ;
        END
        AntennaGateArea 0.1014 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.560 -0.210 7.000 0.210 ;
        RECT  6.300 -0.210 6.560 0.300 ;
        RECT  4.545 -0.210 6.300 0.210 ;
        RECT  4.285 -0.210 4.545 0.300 ;
        RECT  2.750 -0.210 4.285 0.210 ;
        RECT  2.490 -0.210 2.750 0.290 ;
        RECT  2.085 -0.210 2.490 0.210 ;
        RECT  1.825 -0.210 2.085 0.290 ;
        RECT  0.270 -0.210 1.825 0.210 ;
        RECT  0.100 -0.210 0.270 0.745 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.570 2.310 7.000 2.730 ;
        RECT  6.310 2.220 6.570 2.730 ;
        RECT  4.565 2.310 6.310 2.730 ;
        RECT  4.305 2.220 4.565 2.730 ;
        RECT  2.895 2.310 4.305 2.730 ;
        RECT  2.635 2.220 2.895 2.730 ;
        RECT  2.175 2.310 2.635 2.730 ;
        RECT  1.915 2.220 2.175 2.730 ;
        RECT  0.270 2.310 1.915 2.730 ;
        RECT  0.100 1.440 0.270 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.575 0.930 6.670 1.190 ;
        RECT  6.455 0.420 6.575 1.190 ;
        RECT  5.720 0.420 6.455 0.540 ;
        RECT  5.960 0.660 6.150 0.780 ;
        RECT  5.840 0.660 5.960 1.860 ;
        RECT  1.085 1.740 5.840 1.860 ;
        RECT  5.600 0.420 5.720 1.620 ;
        RECT  5.480 1.360 5.600 1.620 ;
        RECT  5.240 0.420 5.360 1.620 ;
        RECT  3.775 0.420 5.240 0.540 ;
        RECT  5.120 1.360 5.240 1.620 ;
        RECT  5.000 0.910 5.120 1.170 ;
        RECT  4.880 0.710 5.000 1.420 ;
        RECT  4.685 0.710 4.880 0.830 ;
        RECT  4.875 1.300 4.880 1.420 ;
        RECT  4.755 1.300 4.875 1.620 ;
        RECT  4.085 1.360 4.205 1.620 ;
        RECT  4.015 0.660 4.155 0.780 ;
        RECT  4.015 1.360 4.085 1.480 ;
        RECT  3.895 0.660 4.015 1.480 ;
        RECT  3.655 0.420 3.775 1.620 ;
        RECT  3.605 0.420 3.655 0.760 ;
        RECT  3.435 0.880 3.535 1.620 ;
        RECT  3.415 0.665 3.435 1.620 ;
        RECT  3.315 0.665 3.415 1.000 ;
        RECT  3.025 1.500 3.415 1.620 ;
        RECT  2.915 0.665 3.315 0.785 ;
        RECT  3.175 1.120 3.295 1.380 ;
        RECT  2.895 1.260 3.175 1.380 ;
        RECT  2.775 1.260 2.895 1.620 ;
        RECT  2.130 1.500 2.775 1.620 ;
        RECT  2.275 0.650 2.395 0.920 ;
        RECT  2.130 0.800 2.275 0.920 ;
        RECT  2.010 0.800 2.130 1.620 ;
        RECT  1.630 1.260 2.010 1.380 ;
        RECT  1.460 1.195 1.630 1.380 ;
        RECT  1.340 1.500 1.630 1.620 ;
        RECT  1.340 0.620 1.495 0.790 ;
        RECT  1.220 0.620 1.340 1.620 ;
        RECT  0.965 0.620 1.085 1.860 ;
        RECT  0.485 0.545 0.605 1.790 ;
    END
END MX4X1AD
MACRO MX4X2AD
    CLASS CORE ;
    FOREIGN MX4X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.195 0.375 7.210 1.645 ;
        RECT  7.050 0.375 7.195 2.005 ;
        RECT  7.025 1.575 7.050 2.005 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.530 1.145 6.650 2.100 ;
        RECT  6.510 1.145 6.530 1.375 ;
        RECT  5.110 1.980 6.530 2.100 ;
        RECT  6.390 1.010 6.510 1.375 ;
        END
        AntennaGateArea 0.2213 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 1.980 4.100 2.100 ;
        RECT  3.390 0.330 3.650 0.545 ;
        RECT  2.940 0.425 3.390 0.545 ;
        RECT  2.820 0.425 2.940 1.140 ;
        RECT  1.920 0.425 2.820 0.545 ;
        RECT  2.350 1.020 2.820 1.140 ;
        RECT  1.800 0.380 1.920 0.545 ;
        RECT  1.730 0.380 1.800 0.500 ;
        RECT  1.470 0.330 1.730 0.500 ;
        RECT  0.860 0.380 1.470 0.500 ;
        RECT  0.740 0.380 0.860 2.170 ;
        RECT  0.585 2.030 0.740 2.170 ;
        END
        AntennaGateArea 0.4364 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 1.110 1.990 1.375 ;
        END
        AntennaGateArea 0.1613 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.100 0.865 0.370 1.290 ;
        RECT  0.070 0.865 0.100 1.095 ;
        END
        AntennaGateArea 0.162 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.105 0.865 3.365 1.140 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.540 0.980 4.790 1.375 ;
        END
        AntennaGateArea 0.161 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.850 -0.210 7.280 0.210 ;
        RECT  6.590 -0.210 6.850 0.390 ;
        RECT  4.990 -0.210 6.590 0.210 ;
        RECT  4.730 -0.210 4.990 0.300 ;
        RECT  3.025 -0.210 4.730 0.210 ;
        RECT  2.765 -0.210 3.025 0.300 ;
        RECT  2.320 -0.210 2.765 0.210 ;
        RECT  2.060 -0.210 2.320 0.305 ;
        RECT  0.295 -0.210 2.060 0.210 ;
        RECT  0.115 -0.210 0.295 0.695 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.810 2.310 7.280 2.730 ;
        RECT  6.550 2.220 6.810 2.730 ;
        RECT  5.110 2.310 6.550 2.730 ;
        RECT  4.850 2.220 5.110 2.730 ;
        RECT  3.090 2.310 4.850 2.730 ;
        RECT  2.830 2.220 3.090 2.730 ;
        RECT  2.325 2.310 2.830 2.730 ;
        RECT  2.065 2.220 2.325 2.730 ;
        RECT  0.310 2.310 2.065 2.730 ;
        RECT  0.130 1.550 0.310 2.730 ;
        RECT  0.000 2.310 0.130 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.280 2.520 ;
        LAYER M1 ;
        RECT  6.810 0.510 6.930 1.240 ;
        RECT  6.155 0.510 6.810 0.630 ;
        RECT  6.270 0.750 6.580 0.870 ;
        RECT  6.270 1.600 6.380 1.860 ;
        RECT  6.150 0.750 6.270 1.860 ;
        RECT  6.000 0.435 6.155 0.630 ;
        RECT  4.860 1.740 6.150 1.860 ;
        RECT  5.880 0.435 6.000 1.620 ;
        RECT  5.640 0.390 5.760 1.575 ;
        RECT  4.140 0.420 5.640 0.540 ;
        RECT  5.495 1.405 5.640 1.575 ;
        RECT  5.325 0.970 5.510 1.230 ;
        RECT  5.060 0.660 5.325 1.620 ;
        RECT  4.740 1.740 4.860 2.100 ;
        RECT  4.370 1.980 4.740 2.100 ;
        RECT  4.490 1.500 4.610 1.860 ;
        RECT  4.380 0.680 4.560 0.800 ;
        RECT  4.380 1.500 4.490 1.620 ;
        RECT  4.260 0.680 4.380 1.620 ;
        RECT  4.250 1.740 4.370 2.100 ;
        RECT  1.100 1.740 4.250 1.860 ;
        RECT  4.130 0.420 4.140 1.620 ;
        RECT  4.010 0.340 4.130 1.620 ;
        RECT  3.770 0.665 3.890 1.620 ;
        RECT  3.495 0.665 3.770 0.835 ;
        RECT  3.260 1.500 3.770 1.620 ;
        RECT  3.515 1.040 3.635 1.380 ;
        RECT  2.660 1.260 3.515 1.380 ;
        RECT  2.230 0.680 2.700 0.800 ;
        RECT  2.490 1.260 2.660 1.575 ;
        RECT  2.230 1.260 2.490 1.380 ;
        RECT  2.110 0.680 2.230 1.380 ;
        RECT  1.610 0.870 2.110 0.990 ;
        RECT  1.340 1.495 1.895 1.615 ;
        RECT  1.340 0.630 1.680 0.750 ;
        RECT  1.490 0.870 1.610 1.300 ;
        RECT  1.220 0.630 1.340 1.615 ;
        RECT  0.980 0.630 1.100 1.860 ;
        RECT  0.500 0.340 0.620 1.910 ;
    END
END MX4X2AD
MACRO MX4X4AD
    CLASS CORE ;
    FOREIGN MX4X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.630 0.805 7.770 1.515 ;
        RECT  7.335 0.805 7.630 0.925 ;
        RECT  7.345 1.395 7.630 1.515 ;
        RECT  7.175 1.395 7.345 2.135 ;
        RECT  7.165 0.420 7.335 0.925 ;
        END
        AntennaDiffArea 0.438 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.530 1.145 6.650 2.100 ;
        RECT  6.510 1.145 6.530 1.375 ;
        RECT  5.110 1.980 6.530 2.100 ;
        RECT  6.390 1.010 6.510 1.375 ;
        END
        AntennaGateArea 0.2213 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 1.980 4.100 2.100 ;
        RECT  3.390 0.330 3.650 0.545 ;
        RECT  2.940 0.425 3.390 0.545 ;
        RECT  2.820 0.425 2.940 1.140 ;
        RECT  1.920 0.425 2.820 0.545 ;
        RECT  2.350 1.020 2.820 1.140 ;
        RECT  1.800 0.380 1.920 0.545 ;
        RECT  1.730 0.380 1.800 0.500 ;
        RECT  1.470 0.330 1.730 0.500 ;
        RECT  0.860 0.380 1.470 0.500 ;
        RECT  0.740 0.380 0.860 2.170 ;
        RECT  0.585 2.030 0.740 2.170 ;
        END
        AntennaGateArea 0.4364 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 1.110 1.990 1.375 ;
        END
        AntennaGateArea 0.1613 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.100 0.865 0.370 1.290 ;
        RECT  0.070 0.865 0.100 1.095 ;
        END
        AntennaGateArea 0.162 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.105 0.865 3.365 1.140 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.540 0.980 4.790 1.375 ;
        END
        AntennaGateArea 0.161 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.705 -0.210 7.840 0.210 ;
        RECT  7.535 -0.210 7.705 0.675 ;
        RECT  7.020 -0.210 7.535 0.210 ;
        RECT  6.760 -0.210 7.020 0.390 ;
        RECT  4.990 -0.210 6.760 0.210 ;
        RECT  4.730 -0.210 4.990 0.300 ;
        RECT  3.025 -0.210 4.730 0.210 ;
        RECT  2.765 -0.210 3.025 0.300 ;
        RECT  2.320 -0.210 2.765 0.210 ;
        RECT  2.060 -0.210 2.320 0.305 ;
        RECT  0.295 -0.210 2.060 0.210 ;
        RECT  0.115 -0.210 0.295 0.695 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.705 2.310 7.840 2.730 ;
        RECT  7.535 1.740 7.705 2.730 ;
        RECT  6.950 2.310 7.535 2.730 ;
        RECT  6.830 1.420 6.950 2.730 ;
        RECT  5.110 2.310 6.830 2.730 ;
        RECT  4.850 2.220 5.110 2.730 ;
        RECT  3.090 2.310 4.850 2.730 ;
        RECT  2.830 2.220 3.090 2.730 ;
        RECT  2.325 2.310 2.830 2.730 ;
        RECT  2.065 2.220 2.325 2.730 ;
        RECT  0.310 2.310 2.065 2.730 ;
        RECT  0.130 1.550 0.310 2.730 ;
        RECT  0.000 2.310 0.130 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.840 2.520 ;
        LAYER M1 ;
        RECT  7.045 1.045 7.465 1.215 ;
        RECT  6.925 0.510 7.045 1.240 ;
        RECT  6.155 0.510 6.925 0.630 ;
        RECT  6.270 0.750 6.580 0.870 ;
        RECT  6.270 1.600 6.380 1.860 ;
        RECT  6.150 0.750 6.270 1.860 ;
        RECT  6.000 0.435 6.155 0.630 ;
        RECT  4.860 1.740 6.150 1.860 ;
        RECT  5.880 0.435 6.000 1.620 ;
        RECT  5.640 0.390 5.760 1.575 ;
        RECT  4.140 0.420 5.640 0.540 ;
        RECT  5.495 1.405 5.640 1.575 ;
        RECT  5.325 0.970 5.510 1.230 ;
        RECT  5.060 0.660 5.325 1.620 ;
        RECT  4.740 1.740 4.860 2.100 ;
        RECT  4.370 1.980 4.740 2.100 ;
        RECT  4.490 1.500 4.610 1.860 ;
        RECT  4.380 0.680 4.560 0.800 ;
        RECT  4.380 1.500 4.490 1.620 ;
        RECT  4.260 0.680 4.380 1.620 ;
        RECT  4.250 1.740 4.370 2.100 ;
        RECT  1.100 1.740 4.250 1.860 ;
        RECT  4.010 0.340 4.140 1.620 ;
        RECT  3.770 0.665 3.890 1.620 ;
        RECT  3.495 0.665 3.770 0.835 ;
        RECT  3.260 1.500 3.770 1.620 ;
        RECT  3.515 1.040 3.635 1.380 ;
        RECT  2.660 1.260 3.515 1.380 ;
        RECT  2.230 0.680 2.700 0.800 ;
        RECT  2.490 1.260 2.660 1.575 ;
        RECT  2.230 1.260 2.490 1.380 ;
        RECT  2.110 0.680 2.230 1.380 ;
        RECT  1.610 0.870 2.110 0.990 ;
        RECT  1.340 1.495 1.895 1.615 ;
        RECT  1.340 0.630 1.680 0.750 ;
        RECT  1.490 0.870 1.610 1.300 ;
        RECT  1.220 0.630 1.340 1.615 ;
        RECT  0.980 0.630 1.100 1.860 ;
        RECT  0.500 0.340 0.620 1.910 ;
    END
END MX4X4AD
MACRO MX4XLAD
    CLASS CORE ;
    FOREIGN MX4XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.530 0.565 6.650 1.680 ;
        RECT  6.490 0.565 6.530 0.825 ;
        RECT  6.465 1.420 6.530 1.680 ;
        END
        AntennaDiffArea 0.146 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.090 1.140 6.155 2.100 ;
        RECT  6.035 0.865 6.090 2.100 ;
        RECT  5.920 0.865 6.035 1.260 ;
        RECT  5.245 1.980 6.035 2.100 ;
        RECT  4.725 1.980 5.245 2.140 ;
        END
        AntennaGateArea 0.1209 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.740 2.020 3.975 2.140 ;
        RECT  3.220 0.330 3.290 0.450 ;
        RECT  3.030 0.330 3.220 0.500 ;
        RECT  2.765 0.380 3.030 0.500 ;
        RECT  2.645 0.380 2.765 0.540 ;
        RECT  2.620 1.980 2.740 2.140 ;
        RECT  2.600 0.420 2.645 0.540 ;
        RECT  0.860 1.980 2.620 2.100 ;
        RECT  2.480 0.420 2.600 1.180 ;
        RECT  1.420 0.420 2.480 0.540 ;
        RECT  2.450 1.060 2.480 1.180 ;
        RECT  2.330 1.060 2.450 1.320 ;
        RECT  1.160 0.340 1.420 0.540 ;
        RECT  0.860 0.420 1.160 0.540 ;
        RECT  0.740 0.420 0.860 2.100 ;
        RECT  0.630 1.145 0.740 1.375 ;
        RECT  0.560 1.950 0.740 2.100 ;
        END
        AntennaGateArea 0.2021 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.705 1.140 1.965 1.415 ;
        END
        AntennaGateArea 0.0724 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.100 1.040 0.270 1.390 ;
        RECT  0.070 1.145 0.100 1.390 ;
        END
        AntennaGateArea 0.0724 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.890 0.865 3.010 1.095 ;
        RECT  2.720 0.865 2.890 1.175 ;
        END
        AntennaGateArea 0.0724 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.100 1.050 4.410 1.375 ;
        END
        AntennaGateArea 0.0724 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.280 -0.210 6.720 0.210 ;
        RECT  6.020 -0.210 6.280 0.300 ;
        RECT  4.495 -0.210 6.020 0.210 ;
        RECT  4.235 -0.210 4.495 0.300 ;
        RECT  2.510 -0.210 4.235 0.210 ;
        RECT  1.990 -0.210 2.510 0.300 ;
        RECT  0.250 -0.210 1.990 0.210 ;
        RECT  0.090 -0.210 0.250 0.880 ;
        RECT  0.000 -0.210 0.090 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.325 2.310 6.720 2.730 ;
        RECT  6.065 2.220 6.325 2.730 ;
        RECT  4.585 2.310 6.065 2.730 ;
        RECT  4.325 2.220 4.585 2.730 ;
        RECT  2.530 2.310 4.325 2.730 ;
        RECT  2.010 2.220 2.530 2.730 ;
        RECT  0.250 2.310 2.010 2.730 ;
        RECT  0.090 1.510 0.250 2.730 ;
        RECT  0.000 2.310 0.090 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.720 2.520 ;
        LAYER M1 ;
        RECT  6.370 0.945 6.410 1.250 ;
        RECT  6.290 0.420 6.370 1.250 ;
        RECT  6.250 0.420 6.290 1.065 ;
        RECT  5.400 0.420 6.250 0.540 ;
        RECT  5.800 1.380 5.915 1.640 ;
        RECT  5.680 0.660 5.800 1.860 ;
        RECT  4.635 1.740 5.680 1.860 ;
        RECT  5.400 1.360 5.535 1.620 ;
        RECT  5.280 0.420 5.400 1.620 ;
        RECT  5.035 0.420 5.155 1.620 ;
        RECT  4.900 0.420 5.035 0.680 ;
        RECT  4.750 0.960 4.905 1.220 ;
        RECT  4.145 0.420 4.900 0.540 ;
        RECT  4.750 1.500 4.885 1.620 ;
        RECT  4.625 0.670 4.750 1.620 ;
        RECT  4.515 1.740 4.635 1.900 ;
        RECT  4.480 0.670 4.625 0.790 ;
        RECT  2.950 1.780 4.515 1.900 ;
        RECT  3.975 1.540 4.195 1.660 ;
        RECT  4.025 0.380 4.145 0.540 ;
        RECT  3.735 0.380 4.025 0.500 ;
        RECT  3.855 0.650 3.975 1.660 ;
        RECT  3.615 0.380 3.735 1.660 ;
        RECT  3.370 0.575 3.615 0.835 ;
        RECT  3.375 0.955 3.495 1.660 ;
        RECT  3.250 0.955 3.375 1.075 ;
        RECT  3.040 1.540 3.375 1.660 ;
        RECT  3.085 1.195 3.255 1.420 ;
        RECT  3.130 0.625 3.250 1.075 ;
        RECT  2.920 0.625 3.130 0.745 ;
        RECT  2.715 1.300 3.085 1.420 ;
        RECT  2.830 1.740 2.950 1.900 ;
        RECT  1.100 1.740 2.830 1.860 ;
        RECT  2.595 1.300 2.715 1.620 ;
        RECT  2.210 1.500 2.595 1.620 ;
        RECT  2.210 0.660 2.360 0.920 ;
        RECT  2.090 0.660 2.210 1.620 ;
        RECT  1.790 0.660 2.090 0.780 ;
        RECT  1.670 0.660 1.790 1.020 ;
        RECT  1.580 0.900 1.670 1.020 ;
        RECT  1.460 0.900 1.580 1.365 ;
        RECT  1.340 0.660 1.550 0.780 ;
        RECT  1.340 1.500 1.550 1.620 ;
        RECT  1.220 0.660 1.340 1.620 ;
        RECT  0.980 0.665 1.100 1.860 ;
        RECT  0.510 0.645 0.620 0.905 ;
        RECT  0.510 1.495 0.620 1.755 ;
        RECT  0.390 0.645 0.510 1.755 ;
    END
END MX4XLAD
MACRO MXI2DX1AD
    CLASS CORE ;
    FOREIGN MXI2DX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.715 0.630 2.730 1.780 ;
        RECT  2.590 0.630 2.715 2.080 ;
        RECT  2.545 0.630 2.590 0.800 ;
        RECT  2.545 1.650 2.590 2.080 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.965 0.780 1.375 ;
        END
        AntennaGateArea 0.0464 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.910 1.750 1.585 ;
        RECT  1.285 0.910 1.630 1.050 ;
        RECT  1.410 1.465 1.630 1.585 ;
        RECT  1.150 1.465 1.410 1.615 ;
        RECT  1.165 0.385 1.285 1.050 ;
        RECT  0.970 0.385 1.165 0.505 ;
        END
        AntennaDiffArea 0.194 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.670 2.170 1.605 ;
        RECT  1.720 0.670 2.030 0.790 ;
        RECT  1.870 1.485 2.030 1.605 ;
        END
        AntennaDiffArea 0.156 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.380 -0.210 2.800 0.210 ;
        RECT  2.120 -0.210 2.380 0.310 ;
        RECT  0.545 -0.210 2.120 0.210 ;
        RECT  0.375 -0.210 0.545 0.495 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.355 2.310 2.800 2.730 ;
        RECT  2.185 1.975 2.355 2.730 ;
        RECT  0.555 2.310 2.185 2.730 ;
        RECT  0.385 1.985 0.555 2.730 ;
        RECT  0.000 2.310 0.385 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.420 0.975 2.445 1.495 ;
        RECT  2.300 0.430 2.420 1.855 ;
        RECT  1.575 0.430 2.300 0.550 ;
        RECT  1.770 1.735 2.300 1.855 ;
        RECT  1.510 1.705 1.770 1.855 ;
        RECT  1.405 0.430 1.575 0.715 ;
        RECT  1.020 1.205 1.510 1.325 ;
        RECT  0.935 1.740 1.105 2.190 ;
        RECT  0.900 0.725 1.020 1.615 ;
        RECT  0.240 1.740 0.935 1.860 ;
        RECT  0.720 0.725 0.900 0.845 ;
        RECT  0.505 1.495 0.900 1.615 ;
        RECT  0.385 1.020 0.505 1.615 ;
        RECT  0.330 1.020 0.385 1.280 ;
        RECT  0.210 0.700 0.265 0.870 ;
        RECT  0.210 1.365 0.240 1.860 ;
        RECT  0.090 0.700 0.210 1.860 ;
    END
END MXI2DX1AD
MACRO MXI2DX2AD
    CLASS CORE ;
    FOREIGN MXI2DX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.715 0.660 2.730 1.780 ;
        RECT  2.590 0.410 2.715 2.080 ;
        RECT  2.545 0.410 2.590 0.840 ;
        RECT  2.545 1.650 2.590 2.080 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.965 0.780 1.375 ;
        END
        AntennaGateArea 0.0724 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.860 1.750 1.525 ;
        RECT  1.285 0.860 1.630 0.980 ;
        RECT  1.385 1.405 1.630 1.525 ;
        RECT  1.340 1.405 1.385 1.655 ;
        RECT  1.220 1.405 1.340 1.925 ;
        RECT  1.165 0.330 1.285 0.980 ;
        RECT  1.190 1.405 1.220 1.655 ;
        RECT  0.970 0.330 1.165 0.450 ;
        END
        AntennaDiffArea 0.27 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.620 2.170 1.605 ;
        RECT  1.720 0.620 2.030 0.740 ;
        RECT  1.870 1.485 2.030 1.605 ;
        END
        AntennaDiffArea 0.266 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.210 2.800 0.210 ;
        RECT  2.070 -0.210 2.330 0.260 ;
        RECT  0.545 -0.210 2.070 0.210 ;
        RECT  0.375 -0.210 0.545 0.495 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.355 2.310 2.800 2.730 ;
        RECT  2.185 1.975 2.355 2.730 ;
        RECT  0.555 2.310 2.185 2.730 ;
        RECT  0.385 1.985 0.555 2.730 ;
        RECT  0.000 2.310 0.385 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.420 1.020 2.445 1.280 ;
        RECT  2.300 0.380 2.420 1.855 ;
        RECT  1.575 0.380 2.300 0.500 ;
        RECT  1.770 1.735 2.300 1.855 ;
        RECT  1.510 1.705 1.770 1.855 ;
        RECT  1.455 0.380 1.575 0.715 ;
        RECT  1.020 1.120 1.510 1.240 ;
        RECT  1.405 0.545 1.455 0.715 ;
        RECT  0.875 1.740 1.070 2.110 ;
        RECT  0.900 0.725 1.020 1.615 ;
        RECT  0.720 0.725 0.900 0.845 ;
        RECT  0.505 1.495 0.900 1.615 ;
        RECT  0.240 1.740 0.875 1.860 ;
        RECT  0.385 1.020 0.505 1.615 ;
        RECT  0.330 1.020 0.385 1.280 ;
        RECT  0.210 0.735 0.265 0.905 ;
        RECT  0.210 1.365 0.240 1.860 ;
        RECT  0.090 0.735 0.210 1.860 ;
    END
END MXI2DX2AD
MACRO MXI2DX4AD
    CLASS CORE ;
    FOREIGN MXI2DX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.755 0.700 3.850 1.540 ;
        RECT  3.710 0.420 3.755 1.955 ;
        RECT  3.585 0.420 3.710 0.850 ;
        RECT  3.585 1.355 3.710 1.955 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.965 0.865 1.375 ;
        END
        AntennaGateArea 0.1444 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.015 0.820 2.090 1.610 ;
        RECT  1.970 0.620 2.015 1.610 ;
        RECT  1.755 0.620 1.970 0.940 ;
        RECT  1.370 1.470 1.970 1.610 ;
        RECT  1.345 0.820 1.755 0.940 ;
        RECT  1.250 1.470 1.370 1.840 ;
        RECT  1.225 0.330 1.345 0.940 ;
        RECT  1.035 0.330 1.225 0.450 ;
        END
        AntennaDiffArea 0.524 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.575 0.620 2.745 1.630 ;
        RECT  2.455 0.620 2.575 0.740 ;
        END
        AntennaDiffArea 0.338 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.090 -0.210 4.200 0.210 ;
        RECT  3.970 -0.210 4.090 0.890 ;
        RECT  3.395 -0.210 3.970 0.210 ;
        RECT  3.225 -0.210 3.395 0.890 ;
        RECT  0.615 -0.210 3.225 0.210 ;
        RECT  0.445 -0.210 0.615 0.745 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.115 2.310 4.200 2.730 ;
        RECT  3.945 1.625 4.115 2.730 ;
        RECT  3.395 2.310 3.945 2.730 ;
        RECT  3.225 2.060 3.395 2.730 ;
        RECT  0.595 2.310 3.225 2.730 ;
        RECT  0.425 2.205 0.595 2.730 ;
        RECT  0.000 2.310 0.425 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  3.005 1.045 3.585 1.215 ;
        RECT  3.005 1.460 3.105 1.920 ;
        RECT  2.885 0.380 3.005 1.920 ;
        RECT  2.285 0.380 2.885 0.500 ;
        RECT  1.585 1.750 2.885 1.920 ;
        RECT  2.165 0.380 2.285 0.670 ;
        RECT  1.585 0.380 2.165 0.500 ;
        RECT  1.105 1.120 1.635 1.290 ;
        RECT  1.465 0.380 1.585 0.680 ;
        RECT  1.060 2.030 1.210 2.150 ;
        RECT  0.985 0.670 1.105 1.615 ;
        RECT  0.940 1.740 1.060 2.150 ;
        RECT  0.760 0.670 0.985 0.790 ;
        RECT  0.470 1.495 0.985 1.615 ;
        RECT  0.230 1.740 0.940 1.860 ;
        RECT  0.350 0.980 0.470 1.615 ;
        RECT  0.110 0.515 0.230 1.860 ;
    END
END MXI2DX4AD
MACRO MXI2DXLAD
    CLASS CORE ;
    FOREIGN MXI2DXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.690 2.730 2.075 ;
        RECT  2.545 0.690 2.590 0.860 ;
        RECT  2.545 1.905 2.590 2.075 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.965 0.780 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.910 1.750 1.540 ;
        RECT  1.285 0.910 1.630 1.050 ;
        RECT  1.340 1.420 1.630 1.540 ;
        RECT  1.220 1.420 1.340 1.810 ;
        RECT  1.165 0.385 1.285 1.050 ;
        RECT  0.980 0.385 1.165 0.505 ;
        END
        AntennaDiffArea 0.151 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.645 2.170 1.725 ;
        RECT  1.720 0.645 2.030 0.765 ;
        RECT  1.870 1.605 2.030 1.725 ;
        END
        AntennaDiffArea 0.114 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.380 -0.210 2.800 0.210 ;
        RECT  2.120 -0.210 2.380 0.285 ;
        RECT  0.545 -0.210 2.120 0.210 ;
        RECT  0.375 -0.210 0.545 0.495 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.400 2.310 2.800 2.730 ;
        RECT  2.140 2.085 2.400 2.730 ;
        RECT  0.555 2.310 2.140 2.730 ;
        RECT  0.385 1.985 0.555 2.730 ;
        RECT  0.000 2.310 0.385 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.420 1.075 2.445 1.595 ;
        RECT  2.300 0.405 2.420 1.965 ;
        RECT  1.575 0.405 2.300 0.525 ;
        RECT  1.725 1.845 2.300 1.965 ;
        RECT  1.555 1.660 1.725 1.965 ;
        RECT  1.455 0.405 1.575 0.790 ;
        RECT  1.020 1.180 1.510 1.300 ;
        RECT  1.405 0.620 1.455 0.790 ;
        RECT  0.840 1.740 1.100 2.190 ;
        RECT  0.900 0.725 1.020 1.615 ;
        RECT  0.720 0.725 0.900 0.845 ;
        RECT  0.505 1.495 0.900 1.615 ;
        RECT  0.240 1.740 0.840 1.860 ;
        RECT  0.385 1.020 0.505 1.615 ;
        RECT  0.330 1.020 0.385 1.280 ;
        RECT  0.210 0.700 0.265 0.870 ;
        RECT  0.210 1.425 0.240 1.860 ;
        RECT  0.090 0.700 0.210 1.860 ;
    END
END MXI2DXLAD
MACRO MXI2X1AD
    CLASS CORE ;
    FOREIGN MXI2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.510 1.740 1.655 1.890 ;
        RECT  1.390 0.415 1.510 1.890 ;
        RECT  1.160 0.415 1.390 0.535 ;
        RECT  1.110 1.740 1.390 1.890 ;
        END
        AntennaDiffArea 0.27 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 2.010 1.610 2.185 ;
        RECT  0.830 2.010 1.350 2.130 ;
        RECT  0.710 1.750 0.830 2.130 ;
        RECT  0.215 1.750 0.710 1.980 ;
        END
        AntennaGateArea 0.1384 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.135 0.770 1.375 ;
        END
        AntennaGateArea 0.0904 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.010 2.170 1.375 ;
        RECT  1.870 1.010 2.030 1.180 ;
        END
        AntennaGateArea 0.09 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.155 -0.210 2.240 0.210 ;
        RECT  1.985 -0.210 2.155 0.775 ;
        RECT  0.670 -0.210 1.985 0.210 ;
        RECT  0.410 -0.210 0.670 0.775 ;
        RECT  0.000 -0.210 0.410 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.135 2.310 2.240 2.730 ;
        RECT  1.965 1.500 2.135 2.730 ;
        RECT  0.585 2.310 1.965 2.730 ;
        RECT  0.415 2.140 0.585 2.730 ;
        RECT  0.000 2.310 0.415 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.750 0.575 1.770 0.835 ;
        RECT  1.630 0.575 1.750 1.620 ;
        RECT  1.150 0.655 1.270 1.615 ;
        RECT  0.985 0.655 1.150 0.775 ;
        RECT  0.750 1.495 1.150 1.615 ;
        RECT  0.910 0.895 1.030 1.325 ;
        RECT  0.815 0.540 0.985 0.775 ;
        RECT  0.240 0.895 0.910 1.015 ;
        RECT  0.190 1.460 0.265 1.630 ;
        RECT  0.190 0.575 0.240 1.015 ;
        RECT  0.070 0.575 0.190 1.630 ;
    END
END MXI2X1AD
MACRO MXI2X2AD
    CLASS CORE ;
    FOREIGN MXI2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.645 2.195 2.075 ;
        RECT  2.025 0.470 2.120 2.075 ;
        RECT  2.000 0.470 2.025 1.910 ;
        RECT  1.405 0.470 2.000 0.640 ;
        RECT  1.500 1.790 2.000 1.910 ;
        RECT  1.380 1.620 1.500 1.910 ;
        RECT  1.240 1.620 1.380 1.740 ;
        END
        AntennaDiffArea 0.842 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.985 2.030 1.350 2.170 ;
        RECT  0.865 1.750 0.985 2.170 ;
        RECT  0.365 1.750 0.865 1.870 ;
        RECT  0.195 1.750 0.365 2.035 ;
        END
        AntennaGateArea 0.2252 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.565 1.085 0.735 1.305 ;
        RECT  0.490 1.145 0.565 1.305 ;
        RECT  0.350 1.145 0.490 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 1.045 3.010 1.375 ;
        RECT  2.530 1.045 2.870 1.215 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.820 -0.210 3.080 0.210 ;
        RECT  2.650 -0.210 2.820 0.785 ;
        RECT  0.670 -0.210 2.650 0.210 ;
        RECT  0.500 -0.210 0.670 0.675 ;
        RECT  0.000 -0.210 0.500 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.915 2.310 3.080 2.730 ;
        RECT  2.745 1.520 2.915 2.730 ;
        RECT  0.670 2.310 2.745 2.730 ;
        RECT  0.500 2.060 0.670 2.730 ;
        RECT  0.000 2.310 0.500 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  2.410 1.405 2.555 2.010 ;
        RECT  2.385 0.415 2.410 2.010 ;
        RECT  2.240 0.415 2.385 1.525 ;
        RECT  1.760 0.760 1.880 1.670 ;
        RECT  1.215 0.760 1.760 0.880 ;
        RECT  1.645 1.380 1.760 1.670 ;
        RECT  1.075 1.380 1.645 1.500 ;
        RECT  1.520 1.000 1.640 1.260 ;
        RECT  0.975 1.000 1.520 1.120 ;
        RECT  1.095 0.590 1.215 0.880 ;
        RECT  1.075 0.590 1.095 0.710 ;
        RECT  0.815 0.330 1.075 0.710 ;
        RECT  0.920 1.380 1.075 1.595 ;
        RECT  0.855 0.830 0.975 1.120 ;
        RECT  0.815 1.475 0.920 1.595 ;
        RECT  0.230 0.830 0.855 0.950 ;
        RECT  0.110 0.640 0.230 1.600 ;
    END
END MXI2X2AD
MACRO MXI2X3AD
    CLASS CORE ;
    FOREIGN MXI2X3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.190 0.670 3.335 1.330 ;
        RECT  3.190 1.535 3.280 1.655 ;
        RECT  3.165 0.670 3.190 1.655 ;
        RECT  3.020 1.160 3.165 1.655 ;
        RECT  2.615 1.160 3.020 1.330 ;
        RECT  2.515 0.415 2.615 1.330 ;
        RECT  2.445 0.415 2.515 1.900 ;
        RECT  1.855 0.415 2.445 0.535 ;
        RECT  2.310 1.160 2.445 1.900 ;
        RECT  1.795 1.780 2.310 1.900 ;
        RECT  1.685 0.415 1.855 0.710 ;
        RECT  1.675 1.610 1.795 1.900 ;
        RECT  1.565 1.610 1.675 1.780 ;
        END
        AntennaDiffArea 0.87 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 2.020 3.530 2.140 ;
        RECT  1.435 1.900 1.555 2.140 ;
        RECT  0.315 1.900 1.435 2.020 ;
        RECT  0.210 1.900 0.315 2.185 ;
        RECT  0.145 1.705 0.210 2.185 ;
        RECT  0.070 1.705 0.145 2.020 ;
        END
        AntennaGateArea 0.3418 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.775 1.085 0.945 1.255 ;
        RECT  0.490 1.085 0.775 1.225 ;
        RECT  0.350 0.865 0.490 1.225 ;
        END
        AntennaGateArea 0.2448 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.895 1.055 4.075 1.175 ;
        RECT  3.555 0.910 3.895 1.175 ;
        END
        AntennaGateArea 0.244 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.080 -0.210 4.480 0.210 ;
        RECT  3.820 -0.210 4.080 0.550 ;
        RECT  1.335 -0.210 3.820 0.210 ;
        RECT  1.165 -0.210 1.335 0.710 ;
        RECT  0.615 -0.210 1.165 0.210 ;
        RECT  0.445 -0.210 0.615 0.745 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.035 2.310 4.480 2.730 ;
        RECT  3.865 1.595 4.035 2.730 ;
        RECT  1.315 2.310 3.865 2.730 ;
        RECT  1.195 2.160 1.315 2.730 ;
        RECT  0.555 2.310 1.195 2.730 ;
        RECT  0.435 2.160 0.555 2.730 ;
        RECT  0.000 2.310 0.435 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
        LAYER M1 ;
        RECT  4.225 0.440 4.395 1.935 ;
        RECT  3.675 0.670 4.225 0.790 ;
        RECT  3.675 1.295 4.225 1.415 ;
        RECT  3.505 0.395 3.675 0.790 ;
        RECT  3.505 1.295 3.675 1.900 ;
        RECT  2.975 0.395 3.505 0.515 ;
        RECT  2.875 1.780 3.505 1.900 ;
        RECT  2.805 0.395 2.975 0.930 ;
        RECT  2.705 1.625 2.875 1.900 ;
        RECT  2.180 0.665 2.215 0.950 ;
        RECT  2.060 0.665 2.180 1.660 ;
        RECT  2.045 0.665 2.060 0.950 ;
        RECT  1.920 1.370 2.060 1.660 ;
        RECT  0.975 0.830 2.045 0.950 ;
        RECT  1.440 1.370 1.920 1.490 ;
        RECT  1.190 1.105 1.670 1.225 ;
        RECT  1.320 1.370 1.440 1.770 ;
        RECT  0.745 1.650 1.320 1.770 ;
        RECT  1.070 1.105 1.190 1.530 ;
        RECT  0.255 1.410 1.070 1.530 ;
        RECT  0.805 0.615 0.975 0.950 ;
        RECT  0.205 0.610 0.255 0.780 ;
        RECT  0.205 1.410 0.255 1.580 ;
        RECT  0.085 0.610 0.205 1.580 ;
    END
END MXI2X3AD
MACRO MXI2X4AD
    CLASS CORE ;
    FOREIGN MXI2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.270 0.860 3.360 0.980 ;
        RECT  3.145 0.860 3.270 1.330 ;
        RECT  3.100 0.860 3.145 1.655 ;
        RECT  2.885 1.160 3.100 1.655 ;
        RECT  2.575 1.160 2.885 1.330 ;
        RECT  2.450 0.620 2.575 1.330 ;
        RECT  2.405 0.620 2.450 1.900 ;
        RECT  1.620 0.620 2.405 0.740 ;
        RECT  2.210 1.160 2.405 1.900 ;
        RECT  1.565 1.780 2.210 1.900 ;
        RECT  1.445 1.640 1.565 1.900 ;
        END
        AntennaDiffArea 1.112 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 2.020 3.415 2.140 ;
        RECT  0.330 2.020 0.400 2.150 ;
        RECT  0.210 1.935 0.330 2.150 ;
        RECT  0.140 1.705 0.210 2.150 ;
        RECT  0.070 1.705 0.140 2.040 ;
        END
        AntennaGateArea 0.4176 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.110 0.835 1.230 ;
        RECT  0.350 0.865 0.490 1.230 ;
        END
        AntennaGateArea 0.3217 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.895 1.055 4.075 1.175 ;
        RECT  3.555 0.910 3.895 1.175 ;
        END
        AntennaGateArea 0.314 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.080 -0.210 4.480 0.210 ;
        RECT  3.820 -0.210 4.080 0.465 ;
        RECT  1.450 -0.210 3.820 0.210 ;
        RECT  1.190 -0.210 1.450 0.260 ;
        RECT  0.615 -0.210 1.190 0.210 ;
        RECT  0.445 -0.210 0.615 0.745 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.035 2.310 4.480 2.730 ;
        RECT  3.865 1.595 4.035 2.730 ;
        RECT  1.385 2.310 3.865 2.730 ;
        RECT  1.125 2.260 1.385 2.730 ;
        RECT  0.625 2.310 1.125 2.730 ;
        RECT  0.365 2.290 0.625 2.730 ;
        RECT  0.000 2.310 0.365 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
        LAYER M1 ;
        RECT  4.225 0.440 4.395 2.185 ;
        RECT  3.720 0.670 4.225 0.790 ;
        RECT  3.720 1.295 4.225 1.415 ;
        RECT  3.565 0.620 3.720 0.790 ;
        RECT  3.460 1.295 3.720 1.900 ;
        RECT  2.935 0.620 3.565 0.740 ;
        RECT  3.270 0.330 3.530 0.500 ;
        RECT  2.740 1.780 3.460 1.900 ;
        RECT  1.500 0.380 3.270 0.500 ;
        RECT  2.765 0.620 2.935 0.800 ;
        RECT  2.570 1.625 2.740 1.900 ;
        RECT  2.065 0.860 2.260 0.980 ;
        RECT  2.015 0.860 2.065 1.490 ;
        RECT  1.945 0.860 2.015 1.660 ;
        RECT  1.020 0.860 1.945 0.980 ;
        RECT  1.755 1.370 1.945 1.660 ;
        RECT  1.315 1.370 1.755 1.490 ;
        RECT  1.075 1.105 1.560 1.225 ;
        RECT  1.380 0.380 1.500 0.740 ;
        RECT  1.195 1.370 1.315 1.770 ;
        RECT  0.745 1.650 1.195 1.770 ;
        RECT  0.955 1.105 1.075 1.530 ;
        RECT  0.900 0.640 1.020 0.980 ;
        RECT  0.255 1.410 0.955 1.530 ;
        RECT  0.760 0.640 0.900 0.760 ;
        RECT  0.205 1.410 0.255 1.580 ;
        RECT  0.205 0.425 0.230 0.945 ;
        RECT  0.085 0.425 0.205 1.580 ;
    END
END MXI2X4AD
MACRO MXI2X6AD
    CLASS CORE ;
    FOREIGN MXI2X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.255 1.420 3.305 1.660 ;
        RECT  3.085 0.625 3.255 1.660 ;
        RECT  2.465 0.625 3.085 0.795 ;
        RECT  1.890 1.510 3.085 1.660 ;
        RECT  2.295 0.365 2.465 0.795 ;
        RECT  1.530 0.625 2.295 0.795 ;
        RECT  1.630 1.510 1.890 1.900 ;
        END
        AntennaDiffArea 1.188 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 1.200 2.410 1.320 ;
        RECT  1.890 1.200 2.060 1.390 ;
        RECT  0.770 1.270 1.890 1.390 ;
        RECT  0.630 1.130 0.770 1.390 ;
        END
        AntennaGateArea 0.6504 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.895 1.100 4.350 1.220 ;
        RECT  3.665 0.910 3.895 1.220 ;
        RECT  3.570 1.100 3.665 1.220 ;
        END
        AntennaGateArea 0.486 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.295 1.055 5.605 1.225 ;
        RECT  5.065 1.055 5.295 1.330 ;
        RECT  4.915 1.055 5.065 1.225 ;
        END
        AntennaGateArea 0.486 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.485 -0.210 6.160 0.210 ;
        RECT  5.225 -0.210 5.485 0.390 ;
        RECT  4.730 -0.210 5.225 0.210 ;
        RECT  4.470 -0.210 4.730 0.390 ;
        RECT  3.925 -0.210 4.470 0.210 ;
        RECT  3.755 -0.210 3.925 0.485 ;
        RECT  1.015 -0.210 3.755 0.210 ;
        RECT  0.845 -0.210 1.015 0.325 ;
        RECT  0.255 -0.210 0.845 0.210 ;
        RECT  0.085 -0.210 0.255 0.380 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.540 2.310 6.160 2.730 ;
        RECT  5.280 2.020 5.540 2.730 ;
        RECT  4.820 2.310 5.280 2.730 ;
        RECT  4.560 2.020 4.820 2.730 ;
        RECT  4.030 2.310 4.560 2.730 ;
        RECT  3.910 2.015 4.030 2.730 ;
        RECT  1.145 2.310 3.910 2.730 ;
        RECT  0.975 2.025 1.145 2.730 ;
        RECT  0.335 2.310 0.975 2.730 ;
        RECT  0.165 2.020 0.335 2.730 ;
        RECT  0.000 2.310 0.165 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.970 0.510 6.090 1.875 ;
        RECT  4.305 0.510 5.970 0.630 ;
        RECT  4.415 1.755 5.970 1.875 ;
        RECT  4.780 0.760 5.845 0.880 ;
        RECT  5.710 1.365 5.830 1.625 ;
        RECT  4.780 1.505 5.710 1.625 ;
        RECT  4.610 0.760 4.780 1.625 ;
        RECT  3.545 1.455 4.610 1.625 ;
        RECT  4.245 1.755 4.415 2.185 ;
        RECT  4.135 0.355 4.305 0.785 ;
        RECT  3.785 1.755 4.245 1.875 ;
        RECT  3.545 0.615 4.135 0.785 ;
        RECT  3.665 1.755 3.785 2.140 ;
        RECT  2.730 2.020 3.665 2.140 ;
        RECT  3.375 0.380 3.545 0.825 ;
        RECT  3.425 1.455 3.545 1.900 ;
        RECT  2.225 1.780 3.425 1.900 ;
        RECT  2.610 0.380 3.375 0.500 ;
        RECT  2.865 1.200 2.955 1.320 ;
        RECT  2.695 0.960 2.865 1.320 ;
        RECT  1.020 0.960 2.695 1.080 ;
        RECT  2.055 1.780 2.225 2.140 ;
        RECT  1.385 0.380 2.150 0.500 ;
        RECT  1.485 2.020 2.055 2.140 ;
        RECT  1.315 1.685 1.485 2.140 ;
        RECT  1.215 0.330 1.385 0.760 ;
        RECT  0.220 1.780 1.315 1.900 ;
        RECT  0.220 0.510 1.215 0.630 ;
        RECT  0.900 0.750 1.020 1.080 ;
        RECT  0.510 0.750 0.900 0.870 ;
        RECT  0.510 1.540 0.760 1.660 ;
        RECT  0.390 0.750 0.510 1.660 ;
        RECT  0.100 0.510 0.220 1.900 ;
    END
END MXI2X6AD
MACRO MXI2X8AD
    CLASS CORE ;
    FOREIGN MXI2X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.610 1.490 4.790 1.660 ;
        RECT  4.130 0.620 4.610 1.660 ;
        RECT  1.470 0.620 4.130 0.780 ;
        RECT  2.505 1.490 4.130 1.660 ;
        RECT  2.245 1.490 2.505 1.770 ;
        RECT  1.785 1.490 2.245 1.660 ;
        RECT  1.525 1.490 1.785 1.755 ;
        END
        AntennaDiffArea 1.794 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.250 2.935 1.370 ;
        RECT  0.920 1.160 1.040 1.370 ;
        RECT  0.550 1.160 0.920 1.330 ;
        END
        AntennaGateArea 0.9163 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.415 1.070 6.725 1.190 ;
        RECT  6.185 0.910 6.415 1.190 ;
        RECT  5.685 1.070 6.185 1.190 ;
        END
        AntennaGateArea 0.648 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.535 1.050 8.080 1.220 ;
        RECT  7.305 1.050 7.535 1.330 ;
        RECT  7.130 1.050 7.305 1.220 ;
        END
        AntennaGateArea 0.648 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.520 -0.210 8.680 0.210 ;
        RECT  8.260 -0.210 8.520 0.390 ;
        RECT  7.780 -0.210 8.260 0.210 ;
        RECT  7.520 -0.210 7.780 0.390 ;
        RECT  7.020 -0.210 7.520 0.210 ;
        RECT  6.760 -0.210 7.020 0.390 ;
        RECT  6.210 -0.210 6.760 0.210 ;
        RECT  6.040 -0.210 6.210 0.535 ;
        RECT  5.535 -0.210 6.040 0.210 ;
        RECT  5.275 -0.210 5.535 0.570 ;
        RECT  1.010 -0.210 5.275 0.210 ;
        RECT  0.890 -0.210 1.010 0.380 ;
        RECT  0.255 -0.210 0.890 0.210 ;
        RECT  0.085 -0.210 0.255 0.335 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.570 2.310 8.680 2.730 ;
        RECT  8.450 1.475 8.570 2.730 ;
        RECT  7.780 2.310 8.450 2.730 ;
        RECT  7.520 2.090 7.780 2.730 ;
        RECT  7.020 2.310 7.520 2.730 ;
        RECT  6.760 2.090 7.020 2.730 ;
        RECT  6.255 2.310 6.760 2.730 ;
        RECT  6.085 1.930 6.255 2.730 ;
        RECT  5.510 2.310 6.085 2.730 ;
        RECT  5.390 1.935 5.510 2.730 ;
        RECT  1.015 2.310 5.390 2.730 ;
        RECT  0.845 1.935 1.015 2.730 ;
        RECT  0.295 2.310 0.845 2.730 ;
        RECT  0.125 1.930 0.295 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.680 2.520 ;
        LAYER M1 ;
        RECT  8.330 0.510 8.400 1.220 ;
        RECT  8.280 0.510 8.330 1.970 ;
        RECT  6.595 0.510 8.280 0.630 ;
        RECT  8.210 1.100 8.280 1.970 ;
        RECT  6.615 1.850 8.210 1.970 ;
        RECT  6.995 0.750 8.160 0.870 ;
        RECT  7.970 1.450 8.090 1.710 ;
        RECT  7.355 1.450 7.970 1.570 ;
        RECT  7.185 1.450 7.355 1.715 ;
        RECT  6.995 1.450 7.185 1.570 ;
        RECT  6.875 0.750 6.995 1.570 ;
        RECT  5.030 1.450 6.875 1.570 ;
        RECT  6.445 1.690 6.615 2.120 ;
        RECT  6.425 0.360 6.595 0.790 ;
        RECT  5.895 1.690 6.445 1.810 ;
        RECT  5.850 0.670 6.425 0.790 ;
        RECT  5.725 1.690 5.895 2.120 ;
        RECT  5.680 0.415 5.850 0.845 ;
        RECT  5.270 1.690 5.725 1.810 ;
        RECT  4.925 0.725 5.680 0.845 ;
        RECT  5.150 1.690 5.270 2.140 ;
        RECT  3.390 2.020 5.150 2.140 ;
        RECT  4.910 1.450 5.030 1.900 ;
        RECT  4.755 0.355 4.925 0.845 ;
        RECT  2.845 1.780 4.910 1.900 ;
        RECT  3.270 0.380 4.755 0.500 ;
        RECT  3.485 1.245 3.955 1.365 ;
        RECT  3.365 0.920 3.485 1.365 ;
        RECT  0.720 0.920 3.365 1.040 ;
        RECT  2.675 1.780 2.845 2.140 ;
        RECT  1.325 0.380 2.810 0.500 ;
        RECT  2.145 2.020 2.675 2.140 ;
        RECT  1.885 1.910 2.145 2.140 ;
        RECT  1.380 2.020 1.885 2.140 ;
        RECT  1.210 1.590 1.380 2.140 ;
        RECT  1.155 0.380 1.325 0.685 ;
        RECT  0.190 1.690 1.210 1.810 ;
        RECT  0.190 0.520 1.155 0.640 ;
        RECT  0.430 0.760 0.720 1.040 ;
        RECT  0.430 1.450 0.700 1.570 ;
        RECT  0.310 0.760 0.430 1.570 ;
        RECT  0.070 0.520 0.190 1.810 ;
    END
END MXI2X8AD
MACRO MXI2XLAD
    CLASS CORE ;
    FOREIGN MXI2XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.390 0.415 1.510 1.890 ;
        RECT  1.200 0.415 1.390 0.535 ;
        RECT  1.110 1.735 1.390 1.890 ;
        END
        AntennaDiffArea 0.198 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 2.010 1.610 2.185 ;
        RECT  0.830 2.010 1.350 2.130 ;
        RECT  0.710 1.860 0.830 2.130 ;
        RECT  0.630 1.860 0.710 1.980 ;
        RECT  0.215 1.750 0.630 1.980 ;
        END
        AntennaGateArea 0.1084 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.135 0.770 1.375 ;
        END
        AntennaGateArea 0.0615 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.000 2.170 1.375 ;
        RECT  1.890 1.000 2.030 1.265 ;
        END
        AntennaGateArea 0.06 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.155 -0.210 2.240 0.210 ;
        RECT  1.985 -0.210 2.155 0.775 ;
        RECT  0.670 -0.210 1.985 0.210 ;
        RECT  0.410 -0.210 0.670 0.720 ;
        RECT  0.000 -0.210 0.410 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.135 2.310 2.240 2.730 ;
        RECT  1.965 1.575 2.135 2.730 ;
        RECT  0.585 2.310 1.965 2.730 ;
        RECT  0.415 2.140 0.585 2.730 ;
        RECT  0.000 2.310 0.415 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.630 0.560 1.770 1.780 ;
        RECT  1.150 0.655 1.270 1.615 ;
        RECT  0.985 0.655 1.150 0.775 ;
        RECT  1.010 1.495 1.150 1.615 ;
        RECT  0.910 0.895 1.030 1.325 ;
        RECT  0.750 1.495 1.010 1.655 ;
        RECT  0.815 0.575 0.985 0.775 ;
        RECT  0.240 0.895 0.910 1.015 ;
        RECT  0.190 1.460 0.265 1.630 ;
        RECT  0.190 0.530 0.240 1.015 ;
        RECT  0.070 0.530 0.190 1.630 ;
    END
END MXI2XLAD
MACRO MXI3X1AD
    CLASS CORE ;
    FOREIGN MXI3X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.710 2.525 0.880 ;
        RECT  2.450 1.410 2.525 1.840 ;
        RECT  2.300 0.710 2.450 1.840 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.830 1.170 4.985 1.690 ;
        END
        AntennaGateArea 0.1203 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.705 0.490 1.975 ;
        RECT  0.315 1.855 0.350 1.975 ;
        RECT  0.145 1.855 0.315 2.090 ;
        END
        AntennaGateArea 0.1058 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.725 1.025 3.015 1.375 ;
        END
        AntennaGateArea 0.0484 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.770 1.145 ;
        END
        AntennaGateArea 0.0574 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.685 0.980 1.890 1.375 ;
        END
        AntennaGateArea 0.0584 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.910 -0.210 5.320 0.210 ;
        RECT  4.650 -0.210 4.910 0.810 ;
        RECT  3.305 -0.210 4.650 0.210 ;
        RECT  3.045 -0.210 3.305 0.310 ;
        RECT  2.190 -0.210 3.045 0.210 ;
        RECT  1.930 -0.210 2.190 0.275 ;
        RECT  0.670 -0.210 1.930 0.210 ;
        RECT  0.410 -0.210 0.670 0.745 ;
        RECT  0.000 -0.210 0.410 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.865 2.310 5.320 2.730 ;
        RECT  4.695 1.825 4.865 2.730 ;
        RECT  3.305 2.310 4.695 2.730 ;
        RECT  3.045 2.210 3.305 2.730 ;
        RECT  2.190 2.310 3.045 2.730 ;
        RECT  1.930 2.210 2.190 2.730 ;
        RECT  0.700 2.310 1.930 2.730 ;
        RECT  0.440 2.095 0.700 2.730 ;
        RECT  0.000 2.310 0.440 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.320 2.520 ;
        LAYER M1 ;
        RECT  5.105 0.665 5.225 2.045 ;
        RECT  5.055 0.665 5.105 1.050 ;
        RECT  5.080 1.785 5.105 2.045 ;
        RECT  4.350 0.930 5.055 1.050 ;
        RECT  4.575 1.190 4.675 1.650 ;
        RECT  4.505 1.190 4.575 2.090 ;
        RECT  4.335 0.630 4.505 0.800 ;
        RECT  4.455 1.530 4.505 2.090 ;
        RECT  1.560 1.970 4.455 2.090 ;
        RECT  4.230 0.930 4.350 1.220 ;
        RECT  4.110 0.680 4.335 0.800 ;
        RECT  4.215 1.430 4.335 1.850 ;
        RECT  4.110 1.430 4.215 1.550 ;
        RECT  3.870 0.440 4.170 0.560 ;
        RECT  3.990 0.680 4.110 1.550 ;
        RECT  3.870 1.680 4.000 1.850 ;
        RECT  3.750 0.440 3.870 1.850 ;
        RECT  2.540 0.440 3.750 0.560 ;
        RECT  3.490 0.680 3.630 1.835 ;
        RECT  3.245 0.785 3.365 1.615 ;
        RECT  2.880 0.785 3.245 0.905 ;
        RECT  2.880 1.495 3.245 1.615 ;
        RECT  2.710 0.735 2.880 0.905 ;
        RECT  2.710 1.495 2.880 1.665 ;
        RECT  2.280 0.390 2.540 0.560 ;
        RECT  2.010 0.735 2.130 1.615 ;
        RECT  1.800 0.735 2.010 0.855 ;
        RECT  1.800 1.495 2.010 1.615 ;
        RECT  1.680 0.530 1.800 0.855 ;
        RECT  1.680 1.495 1.800 1.755 ;
        RECT  1.440 0.625 1.560 2.090 ;
        RECT  1.150 0.625 1.440 0.745 ;
        RECT  1.150 1.755 1.440 1.875 ;
        RECT  1.200 0.890 1.320 1.630 ;
        RECT  1.010 0.890 1.200 1.010 ;
        RECT  0.985 1.510 1.200 1.630 ;
        RECT  0.960 1.130 1.080 1.390 ;
        RECT  0.890 0.570 1.010 1.010 ;
        RECT  0.815 1.510 0.985 1.765 ;
        RECT  0.230 1.270 0.960 1.390 ;
        RECT  0.815 0.570 0.890 0.740 ;
        RECT  0.205 0.600 0.265 0.770 ;
        RECT  0.205 1.270 0.230 1.735 ;
        RECT  0.085 0.600 0.205 1.735 ;
    END
END MXI3X1AD
MACRO MXI3X2AD
    CLASS CORE ;
    FOREIGN MXI3X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.710 2.530 0.880 ;
        RECT  2.450 1.390 2.530 1.820 ;
        RECT  2.300 0.710 2.450 1.820 ;
        END
        AntennaDiffArea 0.341 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.095 0.995 5.265 1.655 ;
        RECT  4.380 1.450 5.095 1.570 ;
        END
        AntennaGateArea 0.1749 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.160 1.705 0.330 2.190 ;
        RECT  0.070 1.705 0.160 1.935 ;
        END
        AntennaGateArea 0.1493 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.725 1.025 3.015 1.375 ;
        END
        AntennaGateArea 0.0524 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.770 1.195 ;
        END
        AntennaGateArea 0.103 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.710 0.980 1.915 1.375 ;
        END
        AntennaGateArea 0.1034 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.930 -0.210 5.600 0.210 ;
        RECT  4.670 -0.210 4.930 0.630 ;
        RECT  3.305 -0.210 4.670 0.210 ;
        RECT  4.665 0.510 4.670 0.630 ;
        RECT  3.045 -0.210 3.305 0.290 ;
        RECT  2.140 -0.210 3.045 0.210 ;
        RECT  1.970 -0.210 2.140 0.575 ;
        RECT  0.670 -0.210 1.970 0.210 ;
        RECT  0.410 -0.210 0.670 0.745 ;
        RECT  0.000 -0.210 0.410 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.145 2.310 5.600 2.730 ;
        RECT  4.975 1.810 5.145 2.730 ;
        RECT  3.310 2.310 4.975 2.730 ;
        RECT  3.050 2.245 3.310 2.730 ;
        RECT  2.145 2.310 3.050 2.730 ;
        RECT  1.885 2.245 2.145 2.730 ;
        RECT  0.625 2.310 1.885 2.730 ;
        RECT  0.505 1.560 0.625 2.730 ;
        RECT  0.000 2.310 0.505 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  5.400 0.675 5.520 1.950 ;
        RECT  5.215 0.675 5.400 0.870 ;
        RECT  5.335 1.780 5.400 1.950 ;
        RECT  4.930 0.750 5.215 0.870 ;
        RECT  4.810 0.750 4.930 1.165 ;
        RECT  4.400 1.045 4.810 1.165 ;
        RECT  4.260 1.725 4.795 1.845 ;
        RECT  4.380 2.005 4.640 2.190 ;
        RECT  4.325 0.645 4.495 0.925 ;
        RECT  4.230 1.045 4.400 1.265 ;
        RECT  1.585 2.005 4.380 2.125 ;
        RECT  4.110 0.805 4.325 0.925 ;
        RECT  4.140 1.385 4.260 1.845 ;
        RECT  3.870 0.410 4.150 0.650 ;
        RECT  4.110 1.385 4.140 1.505 ;
        RECT  3.990 0.805 4.110 1.505 ;
        RECT  3.870 1.625 4.020 1.885 ;
        RECT  3.750 0.410 3.870 1.885 ;
        RECT  2.505 0.410 3.750 0.530 ;
        RECT  3.490 0.650 3.630 1.820 ;
        RECT  3.245 0.785 3.365 1.615 ;
        RECT  2.880 0.785 3.245 0.905 ;
        RECT  2.665 1.495 3.245 1.615 ;
        RECT  2.710 0.675 2.880 0.905 ;
        RECT  2.035 0.735 2.155 1.635 ;
        RECT  1.825 0.735 2.035 0.855 ;
        RECT  1.825 1.515 2.035 1.635 ;
        RECT  1.705 0.430 1.825 0.855 ;
        RECT  1.705 1.515 1.825 1.820 ;
        RECT  1.510 0.430 1.705 0.550 ;
        RECT  1.465 0.670 1.585 2.125 ;
        RECT  1.365 0.670 1.465 0.790 ;
        RECT  1.155 1.825 1.465 1.945 ;
        RECT  1.195 0.610 1.365 0.790 ;
        RECT  1.225 0.910 1.345 1.675 ;
        RECT  1.010 0.910 1.225 1.030 ;
        RECT  1.010 1.555 1.225 1.675 ;
        RECT  0.985 1.150 1.105 1.435 ;
        RECT  0.890 0.570 1.010 1.030 ;
        RECT  0.840 1.555 1.010 2.000 ;
        RECT  0.255 1.315 0.985 1.435 ;
        RECT  0.815 0.570 0.890 0.740 ;
        RECT  0.205 1.315 0.255 1.555 ;
        RECT  0.205 0.555 0.230 0.815 ;
        RECT  0.085 0.555 0.205 1.555 ;
    END
END MXI3X2AD
MACRO MXI3X4AD
    CLASS CORE ;
    FOREIGN MXI3X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.210 0.795 6.370 1.600 ;
        RECT  5.990 0.795 6.210 0.935 ;
        RECT  6.010 1.440 6.210 1.600 ;
        RECT  5.850 1.440 6.010 2.040 ;
        RECT  5.850 0.360 5.990 0.935 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.790 0.865 4.970 1.280 ;
        RECT  4.645 1.110 4.790 1.280 ;
        END
        AntennaGateArea 0.2135 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.025 2.170 1.410 ;
        RECT  1.460 1.110 2.000 1.230 ;
        RECT  1.340 0.900 1.460 1.230 ;
        END
        AntennaGateArea 0.1825 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.945 2.800 1.375 ;
        END
        AntennaGateArea 0.0654 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.860 0.585 1.890 0.870 ;
        RECT  1.695 0.585 1.860 0.990 ;
        RECT  1.600 0.870 1.695 0.990 ;
        END
        AntennaGateArea 0.129 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.980 0.230 1.375 ;
        END
        AntennaGateArea 0.129 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.355 -0.210 6.440 0.210 ;
        RECT  6.185 -0.210 6.355 0.675 ;
        RECT  5.680 -0.210 6.185 0.210 ;
        RECT  5.420 -0.210 5.680 0.390 ;
        RECT  5.050 -0.210 5.420 0.210 ;
        RECT  4.790 -0.210 5.050 0.390 ;
        RECT  3.080 -0.210 4.790 0.210 ;
        RECT  2.820 -0.210 3.080 0.515 ;
        RECT  1.935 -0.210 2.820 0.210 ;
        RECT  1.765 -0.210 1.935 0.465 ;
        RECT  0.230 -0.210 1.765 0.210 ;
        RECT  0.110 -0.210 0.230 0.750 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.370 2.310 6.440 2.730 ;
        RECT  6.210 1.745 6.370 2.730 ;
        RECT  5.680 2.310 6.210 2.730 ;
        RECT  5.420 2.130 5.680 2.730 ;
        RECT  4.980 2.310 5.420 2.730 ;
        RECT  4.720 2.210 4.980 2.730 ;
        RECT  3.100 2.310 4.720 2.730 ;
        RECT  2.840 2.130 3.100 2.730 ;
        RECT  2.050 2.310 2.840 2.730 ;
        RECT  1.790 2.130 2.050 2.730 ;
        RECT  0.230 2.310 1.790 2.730 ;
        RECT  0.070 1.510 0.230 2.730 ;
        RECT  0.000 2.310 0.070 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.440 2.520 ;
        LAYER M1 ;
        RECT  5.715 1.065 5.970 1.185 ;
        RECT  5.595 0.520 5.715 1.185 ;
        RECT  5.490 1.355 5.610 2.010 ;
        RECT  4.490 0.520 5.595 0.640 ;
        RECT  5.455 1.355 5.490 1.475 ;
        RECT  5.220 1.890 5.490 2.010 ;
        RECT  5.335 1.040 5.455 1.475 ;
        RECT  5.215 0.760 5.410 0.880 ;
        RECT  5.215 1.600 5.365 1.770 ;
        RECT  5.100 1.890 5.220 2.090 ;
        RECT  5.095 0.760 5.215 1.770 ;
        RECT  4.500 1.970 5.100 2.090 ;
        RECT  4.980 1.650 5.095 1.770 ;
        RECT  4.860 1.650 4.980 1.845 ;
        RECT  3.990 1.725 4.860 1.845 ;
        RECT  4.335 1.485 4.740 1.605 ;
        RECT  4.335 0.760 4.665 0.880 ;
        RECT  4.380 1.970 4.500 2.140 ;
        RECT  4.370 0.380 4.490 0.640 ;
        RECT  3.345 2.020 4.380 2.140 ;
        RECT  3.750 0.380 4.370 0.500 ;
        RECT  4.215 0.760 4.335 1.605 ;
        RECT  3.990 0.620 4.095 0.880 ;
        RECT  3.870 0.620 3.990 1.845 ;
        RECT  3.610 0.380 3.750 1.890 ;
        RECT  3.250 0.360 3.390 1.750 ;
        RECT  3.225 1.890 3.345 2.140 ;
        RECT  0.900 1.890 3.225 2.010 ;
        RECT  3.010 0.635 3.130 1.615 ;
        RECT  2.650 0.635 3.010 0.755 ;
        RECT  2.650 1.495 3.010 1.615 ;
        RECT  2.530 0.395 2.650 0.755 ;
        RECT  2.530 1.495 2.650 1.755 ;
        RECT  2.290 0.565 2.410 1.710 ;
        RECT  2.145 0.565 2.290 0.735 ;
        RECT  0.950 1.590 2.290 1.710 ;
        RECT  1.260 0.350 1.520 0.755 ;
        RECT  1.190 1.350 1.520 1.470 ;
        RECT  1.190 0.610 1.260 0.755 ;
        RECT  1.070 0.610 1.190 1.470 ;
        RECT  0.830 0.465 0.950 0.850 ;
        RECT  0.830 0.980 0.950 1.710 ;
        RECT  0.780 1.830 0.900 2.010 ;
        RECT  0.710 0.730 0.830 0.850 ;
        RECT  0.710 1.830 0.780 1.950 ;
        RECT  0.590 0.730 0.710 1.950 ;
        RECT  0.470 2.070 0.660 2.190 ;
        RECT  0.470 0.435 0.615 0.605 ;
        RECT  0.350 0.435 0.470 2.190 ;
    END
END MXI3X4AD
MACRO MXI3XLAD
    CLASS CORE ;
    FOREIGN MXI3XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.455 1.585 2.560 1.845 ;
        RECT  2.455 0.735 2.525 0.905 ;
        RECT  2.305 0.735 2.455 1.845 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.830 1.145 4.970 1.655 ;
        END
        AntennaGateArea 0.0969 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.705 0.490 2.075 ;
        RECT  0.145 1.905 0.350 2.075 ;
        END
        AntennaGateArea 0.0968 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.145 3.125 1.375 ;
        END
        AntennaGateArea 0.0484 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.770 1.125 ;
        END
        AntennaGateArea 0.0484 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 0.865 1.890 1.390 ;
        END
        AntennaGateArea 0.0484 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.910 -0.210 5.320 0.210 ;
        RECT  4.650 -0.210 4.910 0.785 ;
        RECT  3.320 -0.210 4.650 0.210 ;
        RECT  3.060 -0.210 3.320 0.310 ;
        RECT  2.180 -0.210 3.060 0.210 ;
        RECT  1.920 -0.210 2.180 0.310 ;
        RECT  0.670 -0.210 1.920 0.210 ;
        RECT  0.410 -0.210 0.670 0.725 ;
        RECT  0.000 -0.210 0.410 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.830 2.310 5.320 2.730 ;
        RECT  4.710 1.775 4.830 2.730 ;
        RECT  3.360 2.310 4.710 2.730 ;
        RECT  3.100 2.210 3.360 2.730 ;
        RECT  2.250 2.310 3.100 2.730 ;
        RECT  1.990 2.210 2.250 2.730 ;
        RECT  0.870 2.310 1.990 2.730 ;
        RECT  0.610 2.065 0.870 2.730 ;
        RECT  0.000 2.310 0.610 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.320 2.520 ;
        LAYER M1 ;
        RECT  5.090 0.595 5.210 1.835 ;
        RECT  5.055 0.595 5.090 1.025 ;
        RECT  4.390 0.905 5.055 1.025 ;
        RECT  4.420 1.970 4.590 2.150 ;
        RECT  4.150 0.665 4.530 0.785 ;
        RECT  4.325 1.310 4.445 1.805 ;
        RECT  1.560 1.970 4.420 2.090 ;
        RECT  4.270 0.905 4.390 1.190 ;
        RECT  4.150 1.310 4.325 1.430 ;
        RECT  3.910 0.415 4.150 0.535 ;
        RECT  4.030 0.665 4.150 1.430 ;
        RECT  3.910 1.625 4.110 1.795 ;
        RECT  3.790 0.415 3.910 1.795 ;
        RECT  2.510 0.440 3.790 0.560 ;
        RECT  3.550 0.690 3.670 1.835 ;
        RECT  3.310 0.785 3.430 1.720 ;
        RECT  2.885 0.785 3.310 0.905 ;
        RECT  2.980 1.600 3.310 1.720 ;
        RECT  2.720 1.600 2.980 1.745 ;
        RECT  2.715 0.735 2.885 0.905 ;
        RECT  2.250 0.440 2.510 0.590 ;
        RECT  2.010 0.440 2.130 1.630 ;
        RECT  1.510 0.440 2.010 0.560 ;
        RECT  1.800 1.510 2.010 1.630 ;
        RECT  1.680 1.510 1.800 1.770 ;
        RECT  1.440 0.680 1.560 2.090 ;
        RECT  1.345 0.680 1.440 0.800 ;
        RECT  1.090 1.790 1.440 1.910 ;
        RECT  1.175 0.580 1.345 0.800 ;
        RECT  1.200 0.920 1.320 1.670 ;
        RECT  1.010 0.920 1.200 1.040 ;
        RECT  0.900 1.550 1.200 1.670 ;
        RECT  0.960 1.160 1.080 1.430 ;
        RECT  0.890 0.580 1.010 1.040 ;
        RECT  0.230 1.310 0.960 1.430 ;
        RECT  0.780 1.550 0.900 1.810 ;
        RECT  0.815 0.580 0.890 0.750 ;
        RECT  0.205 0.580 0.265 0.750 ;
        RECT  0.205 1.310 0.230 1.740 ;
        RECT  0.085 0.580 0.205 1.740 ;
    END
END MXI3XLAD
MACRO MXI4X1AD
    CLASS CORE ;
    FOREIGN MXI4X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.770 0.650 6.930 1.920 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.855 1.145 5.935 1.405 ;
        RECT  5.670 1.145 5.855 1.655 ;
        END
        AntennaGateArea 0.1218 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.125 2.170 1.495 ;
        END
        AntennaGateArea 0.1655 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 1.125 2.460 1.490 ;
        END
        AntennaGateArea 0.0574 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.690 0.980 3.850 1.375 ;
        RECT  3.585 0.980 3.690 1.360 ;
        END
        AntennaGateArea 0.0587 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.390 0.865 1.650 1.165 ;
        END
        AntennaGateArea 0.0574 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.160 0.845 0.280 1.365 ;
        RECT  0.070 0.845 0.160 1.095 ;
        END
        AntennaGateArea 0.0574 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.620 -0.210 7.000 0.210 ;
        RECT  6.360 -0.210 6.620 0.285 ;
        RECT  5.730 -0.210 6.360 0.210 ;
        RECT  5.560 -0.210 5.730 0.450 ;
        RECT  3.995 -0.210 5.560 0.210 ;
        RECT  3.735 -0.210 3.995 0.310 ;
        RECT  2.450 -0.210 3.735 0.210 ;
        RECT  2.280 -0.210 2.450 0.765 ;
        RECT  1.770 -0.210 2.280 0.210 ;
        RECT  1.510 -0.210 1.770 0.745 ;
        RECT  0.230 -0.210 1.510 0.210 ;
        RECT  0.070 -0.210 0.230 0.585 ;
        RECT  0.000 -0.210 0.070 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.555 2.310 7.000 2.730 ;
        RECT  6.385 1.400 6.555 2.730 ;
        RECT  5.720 2.310 6.385 2.730 ;
        RECT  5.550 1.775 5.720 2.730 ;
        RECT  3.980 2.310 5.550 2.730 ;
        RECT  3.720 2.210 3.980 2.730 ;
        RECT  2.420 2.310 3.720 2.730 ;
        RECT  2.160 2.095 2.420 2.730 ;
        RECT  1.790 2.310 2.160 2.730 ;
        RECT  1.530 2.095 1.790 2.730 ;
        RECT  0.335 2.310 1.530 2.730 ;
        RECT  0.165 2.100 0.335 2.730 ;
        RECT  0.000 2.310 0.165 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.530 0.405 6.650 1.260 ;
        RECT  5.970 0.405 6.530 0.525 ;
        RECT  6.090 0.650 6.210 1.930 ;
        RECT  5.290 0.810 6.090 0.930 ;
        RECT  6.030 1.760 6.090 1.930 ;
        RECT  5.850 0.405 5.970 0.690 ;
        RECT  5.390 0.570 5.850 0.690 ;
        RECT  5.415 1.055 5.535 1.485 ;
        RECT  5.300 1.365 5.415 1.485 ;
        RECT  5.270 0.380 5.390 0.690 ;
        RECT  5.180 1.365 5.300 2.135 ;
        RECT  5.170 0.810 5.290 1.245 ;
        RECT  4.700 0.380 5.270 0.500 ;
        RECT  4.305 2.015 5.180 2.135 ;
        RECT  5.115 0.985 5.170 1.245 ;
        RECT  4.990 1.565 5.060 1.825 ;
        RECT  4.990 0.620 5.050 0.880 ;
        RECT  4.870 0.620 4.990 1.825 ;
        RECT  4.570 0.380 4.700 1.835 ;
        RECT  4.245 0.560 4.365 1.850 ;
        RECT  4.185 1.970 4.305 2.135 ;
        RECT  4.210 0.560 4.245 0.820 ;
        RECT  4.220 1.590 4.245 1.850 ;
        RECT  2.670 1.970 4.185 2.090 ;
        RECT  4.090 0.965 4.125 1.485 ;
        RECT  3.970 0.430 4.090 1.850 ;
        RECT  3.180 0.430 3.970 0.550 ;
        RECT  3.115 1.730 3.970 1.850 ;
        RECT  3.465 0.670 3.615 0.790 ;
        RECT  3.465 1.490 3.570 1.610 ;
        RECT  3.345 0.670 3.465 1.610 ;
        RECT  3.310 1.490 3.345 1.610 ;
        RECT  3.060 0.430 3.180 0.820 ;
        RECT  3.040 0.940 3.160 1.560 ;
        RECT  2.945 1.680 3.115 1.850 ;
        RECT  2.940 0.940 3.040 1.060 ;
        RECT  2.800 1.440 3.040 1.560 ;
        RECT  2.820 0.640 2.940 1.060 ;
        RECT  2.700 1.200 2.920 1.320 ;
        RECT  2.590 0.640 2.820 0.760 ;
        RECT  2.680 1.440 2.800 1.735 ;
        RECT  2.580 0.885 2.700 1.320 ;
        RECT  2.540 1.615 2.680 1.735 ;
        RECT  2.550 1.855 2.670 2.090 ;
        RECT  2.085 0.885 2.580 1.005 ;
        RECT  1.050 1.855 2.550 1.975 ;
        RECT  1.890 1.615 2.170 1.735 ;
        RECT  1.915 0.600 2.085 1.005 ;
        RECT  1.890 0.885 1.915 1.005 ;
        RECT  1.770 0.885 1.890 1.735 ;
        RECT  1.250 1.285 1.770 1.405 ;
        RECT  1.170 1.525 1.340 1.720 ;
        RECT  1.240 0.340 1.310 0.600 ;
        RECT  1.130 1.105 1.250 1.405 ;
        RECT  1.120 0.340 1.240 0.980 ;
        RECT  1.010 1.525 1.170 1.645 ;
        RECT  1.010 0.860 1.120 0.980 ;
        RECT  0.770 1.765 1.050 1.975 ;
        RECT  0.890 0.860 1.010 1.645 ;
        RECT  0.830 0.350 0.950 0.740 ;
        RECT  0.770 0.620 0.830 0.740 ;
        RECT  0.650 0.620 0.770 1.975 ;
        RECT  0.530 0.380 0.660 0.500 ;
        RECT  0.400 0.380 0.530 1.855 ;
    END
END MXI4X1AD
MACRO MXI4X2AD
    CLASS CORE ;
    FOREIGN MXI4X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.770 0.340 6.930 2.160 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.670 1.100 5.995 1.550 ;
        END
        AntennaGateArea 0.1818 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.090 2.170 1.495 ;
        END
        AntennaGateArea 0.2884 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 1.105 2.460 1.490 ;
        END
        AntennaGateArea 0.1034 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.900 3.850 1.375 ;
        END
        AntennaGateArea 0.1034 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.390 0.865 1.650 1.165 ;
        END
        AntennaGateArea 0.1034 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.160 0.780 0.280 1.300 ;
        RECT  0.070 0.865 0.160 1.095 ;
        END
        AntennaGateArea 0.1034 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.530 -0.210 7.000 0.210 ;
        RECT  6.270 -0.210 6.530 0.330 ;
        RECT  5.780 -0.210 6.270 0.210 ;
        RECT  5.610 -0.210 5.780 0.450 ;
        RECT  3.995 -0.210 5.610 0.210 ;
        RECT  3.735 -0.210 3.995 0.310 ;
        RECT  2.400 -0.210 3.735 0.210 ;
        RECT  2.280 -0.210 2.400 0.710 ;
        RECT  1.770 -0.210 2.280 0.210 ;
        RECT  1.510 -0.210 1.770 0.720 ;
        RECT  0.255 -0.210 1.510 0.210 ;
        RECT  0.095 -0.210 0.255 0.650 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.530 2.310 7.000 2.730 ;
        RECT  6.410 1.450 6.530 2.730 ;
        RECT  5.745 2.310 6.410 2.730 ;
        RECT  5.575 1.695 5.745 2.730 ;
        RECT  4.015 2.310 5.575 2.730 ;
        RECT  3.755 2.260 4.015 2.730 ;
        RECT  2.420 2.310 3.755 2.730 ;
        RECT  2.160 2.095 2.420 2.730 ;
        RECT  1.790 2.310 2.160 2.730 ;
        RECT  1.530 2.140 1.790 2.730 ;
        RECT  0.290 2.310 1.530 2.730 ;
        RECT  0.120 2.205 0.290 2.730 ;
        RECT  0.000 2.310 0.120 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.530 0.450 6.650 1.260 ;
        RECT  6.020 0.450 6.530 0.570 ;
        RECT  6.235 0.690 6.305 0.950 ;
        RECT  6.140 0.690 6.235 1.985 ;
        RECT  6.115 0.830 6.140 1.985 ;
        RECT  5.290 0.830 6.115 0.950 ;
        RECT  6.000 1.815 6.115 1.985 ;
        RECT  5.900 0.450 6.020 0.690 ;
        RECT  5.390 0.570 5.900 0.690 ;
        RECT  5.455 1.090 5.535 1.570 ;
        RECT  5.415 1.090 5.455 2.140 ;
        RECT  5.335 1.450 5.415 2.140 ;
        RECT  5.270 0.430 5.390 0.690 ;
        RECT  2.765 2.020 5.335 2.140 ;
        RECT  5.170 0.830 5.290 1.300 ;
        RECT  4.690 0.430 5.270 0.550 ;
        RECT  5.095 1.590 5.215 1.850 ;
        RECT  5.115 1.040 5.170 1.300 ;
        RECT  4.990 1.590 5.095 1.710 ;
        RECT  4.990 0.670 5.050 0.930 ;
        RECT  4.870 0.670 4.990 1.710 ;
        RECT  4.690 1.600 4.740 1.860 ;
        RECT  4.570 0.430 4.690 1.860 ;
        RECT  4.255 0.440 4.375 1.850 ;
        RECT  4.210 0.440 4.255 0.700 ;
        RECT  4.225 1.590 4.255 1.850 ;
        RECT  4.090 1.120 4.135 1.380 ;
        RECT  3.970 0.430 4.090 1.900 ;
        RECT  3.180 0.430 3.970 0.550 ;
        RECT  2.920 1.780 3.970 1.900 ;
        RECT  3.465 1.540 3.635 1.660 ;
        RECT  3.465 0.670 3.615 0.790 ;
        RECT  3.345 0.670 3.465 1.660 ;
        RECT  3.105 0.900 3.225 1.640 ;
        RECT  3.060 0.430 3.180 0.760 ;
        RECT  2.940 0.900 3.105 1.020 ;
        RECT  2.800 1.520 3.105 1.640 ;
        RECT  2.850 1.140 2.970 1.400 ;
        RECT  2.820 0.610 2.940 1.020 ;
        RECT  2.700 1.140 2.850 1.260 ;
        RECT  2.570 0.610 2.820 0.730 ;
        RECT  2.675 1.520 2.800 1.735 ;
        RECT  2.645 1.855 2.765 2.140 ;
        RECT  2.580 0.850 2.700 1.260 ;
        RECT  2.540 1.615 2.675 1.735 ;
        RECT  1.050 1.855 2.645 1.975 ;
        RECT  2.085 0.850 2.580 0.970 ;
        RECT  1.890 1.615 2.170 1.735 ;
        RECT  1.915 0.610 2.085 0.970 ;
        RECT  1.890 0.850 1.915 0.970 ;
        RECT  1.770 0.850 1.890 1.735 ;
        RECT  1.250 1.285 1.770 1.405 ;
        RECT  1.195 1.525 1.365 1.710 ;
        RECT  1.240 0.470 1.310 0.730 ;
        RECT  1.130 1.105 1.250 1.405 ;
        RECT  1.120 0.470 1.240 0.980 ;
        RECT  1.010 1.525 1.195 1.645 ;
        RECT  1.010 0.860 1.120 0.980 ;
        RECT  0.770 1.765 1.050 1.975 ;
        RECT  0.890 0.860 1.010 1.645 ;
        RECT  0.830 0.350 0.950 0.740 ;
        RECT  0.770 0.620 0.830 0.740 ;
        RECT  0.650 0.620 0.770 1.975 ;
        RECT  0.530 0.380 0.660 0.500 ;
        RECT  0.400 0.380 0.530 1.990 ;
    END
END MXI4X2AD
MACRO MXI4X4AD
    CLASS CORE ;
    FOREIGN MXI4X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.090 0.685 7.210 1.550 ;
        RECT  7.060 0.355 7.090 2.155 ;
        RECT  6.970 0.355 7.060 0.875 ;
        RECT  6.970 1.375 7.060 2.155 ;
        END
        AntennaDiffArea 0.442 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.625 0.910 5.860 1.290 ;
        END
        AntennaGateArea 0.2144 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.070 2.170 1.495 ;
        END
        AntennaGateArea 0.3614 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 1.070 2.460 1.490 ;
        END
        AntennaGateArea 0.1124 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.565 1.030 3.850 1.375 ;
        END
        AntennaGateArea 0.1296 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.390 0.865 1.650 1.190 ;
        END
        AntennaGateArea 0.1124 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.155 0.865 0.280 1.325 ;
        RECT  0.070 0.865 0.155 1.100 ;
        END
        AntennaGateArea 0.1204 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.450 -0.210 7.560 0.210 ;
        RECT  7.330 -0.210 7.450 0.855 ;
        RECT  6.750 -0.210 7.330 0.210 ;
        RECT  6.490 -0.210 6.750 0.390 ;
        RECT  6.030 -0.210 6.490 0.210 ;
        RECT  5.770 -0.210 6.030 0.270 ;
        RECT  3.995 -0.210 5.770 0.210 ;
        RECT  3.735 -0.210 3.995 0.410 ;
        RECT  2.425 -0.210 3.735 0.210 ;
        RECT  2.255 -0.210 2.425 0.665 ;
        RECT  1.770 -0.210 2.255 0.210 ;
        RECT  1.510 -0.210 1.770 0.630 ;
        RECT  0.255 -0.210 1.510 0.210 ;
        RECT  0.095 -0.210 0.255 0.650 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.450 2.310 7.560 2.730 ;
        RECT  7.330 1.445 7.450 2.730 ;
        RECT  6.800 2.310 7.330 2.730 ;
        RECT  6.540 2.130 6.800 2.730 ;
        RECT  5.995 2.310 6.540 2.730 ;
        RECT  5.825 2.130 5.995 2.730 ;
        RECT  3.965 2.310 5.825 2.730 ;
        RECT  3.705 2.260 3.965 2.730 ;
        RECT  2.420 2.310 3.705 2.730 ;
        RECT  2.160 2.095 2.420 2.730 ;
        RECT  1.790 2.310 2.160 2.730 ;
        RECT  1.530 2.140 1.790 2.730 ;
        RECT  0.285 2.310 1.530 2.730 ;
        RECT  0.115 2.265 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  6.830 1.025 6.940 1.195 ;
        RECT  6.710 0.510 6.830 1.195 ;
        RECT  5.950 0.510 6.710 0.630 ;
        RECT  6.560 1.250 6.580 2.010 ;
        RECT  6.460 0.990 6.560 2.010 ;
        RECT  6.440 0.990 6.460 1.370 ;
        RECT  5.665 1.890 6.460 2.010 ;
        RECT  6.300 0.760 6.370 0.880 ;
        RECT  6.300 1.510 6.340 1.770 ;
        RECT  6.180 0.760 6.300 1.770 ;
        RECT  6.110 0.760 6.180 0.880 ;
        RECT  5.330 1.650 6.180 1.770 ;
        RECT  5.795 0.390 5.950 0.630 ;
        RECT  4.705 0.390 5.795 0.510 ;
        RECT  5.330 1.410 5.725 1.530 ;
        RECT  5.545 1.890 5.665 2.140 ;
        RECT  5.330 0.630 5.660 0.750 ;
        RECT  2.765 2.020 5.545 2.140 ;
        RECT  5.210 0.630 5.330 1.530 ;
        RECT  5.160 1.650 5.330 1.875 ;
        RECT  4.975 1.650 5.160 1.770 ;
        RECT  4.975 0.665 5.060 0.925 ;
        RECT  4.855 0.665 4.975 1.770 ;
        RECT  4.570 0.390 4.705 1.860 ;
        RECT  4.255 0.440 4.375 1.850 ;
        RECT  4.210 0.440 4.255 0.700 ;
        RECT  4.225 1.590 4.255 1.850 ;
        RECT  4.090 1.120 4.135 1.380 ;
        RECT  3.970 0.540 4.090 1.900 ;
        RECT  3.180 0.540 3.970 0.660 ;
        RECT  2.920 1.780 3.970 1.900 ;
        RECT  3.360 0.780 3.615 0.900 ;
        RECT  3.360 1.540 3.540 1.660 ;
        RECT  3.240 0.780 3.360 1.660 ;
        RECT  3.060 0.370 3.180 0.660 ;
        RECT  3.000 0.850 3.120 1.640 ;
        RECT  2.940 0.850 3.000 0.970 ;
        RECT  2.800 1.520 3.000 1.640 ;
        RECT  2.820 0.535 2.940 0.970 ;
        RECT  2.760 1.090 2.880 1.350 ;
        RECT  2.785 0.535 2.820 0.655 ;
        RECT  2.675 1.520 2.800 1.735 ;
        RECT  2.615 0.485 2.785 0.655 ;
        RECT  2.645 1.855 2.765 2.140 ;
        RECT  2.700 1.090 2.760 1.210 ;
        RECT  2.580 0.815 2.700 1.210 ;
        RECT  2.540 1.615 2.675 1.735 ;
        RECT  0.770 1.855 2.645 1.975 ;
        RECT  2.085 0.815 2.580 0.935 ;
        RECT  1.890 1.615 2.170 1.735 ;
        RECT  1.915 0.610 2.085 0.935 ;
        RECT  1.890 0.815 1.915 0.935 ;
        RECT  1.770 0.815 1.890 1.735 ;
        RECT  1.250 1.310 1.770 1.430 ;
        RECT  1.010 1.565 1.410 1.685 ;
        RECT  1.240 0.470 1.310 0.730 ;
        RECT  1.130 1.070 1.250 1.430 ;
        RECT  1.120 0.470 1.240 0.935 ;
        RECT  1.010 0.815 1.120 0.935 ;
        RECT  0.890 0.815 1.010 1.685 ;
        RECT  0.830 0.350 0.950 0.695 ;
        RECT  0.770 0.575 0.830 0.695 ;
        RECT  0.650 0.575 0.770 1.975 ;
        RECT  0.530 0.330 0.660 0.450 ;
        RECT  0.400 0.330 0.530 2.010 ;
    END
END MXI4X4AD
MACRO MXI4XLAD
    CLASS CORE ;
    FOREIGN MXI4XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.760 0.690 6.930 1.695 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.855 1.145 5.980 1.405 ;
        RECT  5.670 1.145 5.855 1.655 ;
        END
        AntennaGateArea 0.0976 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.125 2.170 1.495 ;
        END
        AntennaGateArea 0.147 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.125 2.460 1.655 ;
        END
        AntennaGateArea 0.0489 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 0.930 3.850 1.375 ;
        END
        AntennaGateArea 0.0501 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.390 0.865 1.650 1.165 ;
        END
        AntennaGateArea 0.0484 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.170 0.835 0.290 1.355 ;
        RECT  0.070 0.835 0.170 1.095 ;
        END
        AntennaGateArea 0.0484 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.630 -0.210 7.000 0.210 ;
        RECT  6.370 -0.210 6.630 0.285 ;
        RECT  5.730 -0.210 6.370 0.210 ;
        RECT  5.560 -0.210 5.730 0.450 ;
        RECT  4.050 -0.210 5.560 0.210 ;
        RECT  3.790 -0.210 4.050 0.310 ;
        RECT  2.455 -0.210 3.790 0.210 ;
        RECT  2.285 -0.210 2.455 0.765 ;
        RECT  1.735 -0.210 2.285 0.210 ;
        RECT  1.565 -0.210 1.735 0.745 ;
        RECT  0.265 -0.210 1.565 0.210 ;
        RECT  0.095 -0.210 0.265 0.570 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.555 2.310 7.000 2.730 ;
        RECT  6.385 1.435 6.555 2.730 ;
        RECT  5.825 2.310 6.385 2.730 ;
        RECT  5.655 1.775 5.825 2.730 ;
        RECT  4.030 2.310 5.655 2.730 ;
        RECT  3.770 2.210 4.030 2.730 ;
        RECT  2.470 2.310 3.770 2.730 ;
        RECT  2.210 2.095 2.470 2.730 ;
        RECT  1.790 2.310 2.210 2.730 ;
        RECT  1.530 2.095 1.790 2.730 ;
        RECT  0.335 2.310 1.530 2.730 ;
        RECT  0.165 2.060 0.335 2.730 ;
        RECT  0.000 2.310 0.165 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.520 0.405 6.640 1.260 ;
        RECT  5.970 0.405 6.520 0.525 ;
        RECT  6.100 0.650 6.220 1.915 ;
        RECT  5.440 0.905 6.100 1.025 ;
        RECT  6.045 1.745 6.100 1.915 ;
        RECT  5.850 0.405 5.970 0.690 ;
        RECT  5.440 0.570 5.850 0.690 ;
        RECT  2.720 1.970 5.535 2.090 ;
        RECT  5.320 0.380 5.440 0.690 ;
        RECT  5.320 0.905 5.440 1.120 ;
        RECT  4.990 1.640 5.415 1.770 ;
        RECT  4.750 0.380 5.320 0.500 ;
        RECT  5.235 1.000 5.320 1.120 ;
        RECT  5.115 1.000 5.235 1.520 ;
        RECT  5.080 0.620 5.200 0.880 ;
        RECT  4.990 0.760 5.080 0.880 ;
        RECT  4.870 0.760 4.990 1.770 ;
        RECT  4.630 0.380 4.750 1.835 ;
        RECT  4.580 1.575 4.630 1.835 ;
        RECT  4.340 0.575 4.380 0.835 ;
        RECT  4.220 0.575 4.340 1.850 ;
        RECT  3.980 0.430 4.100 1.850 ;
        RECT  3.185 0.430 3.980 0.550 ;
        RECT  3.230 1.730 3.980 1.850 ;
        RECT  3.480 1.490 3.620 1.610 ;
        RECT  3.480 0.670 3.590 0.840 ;
        RECT  3.360 0.670 3.480 1.610 ;
        RECT  2.970 1.685 3.230 1.850 ;
        RECT  3.090 0.960 3.210 1.560 ;
        RECT  3.065 0.430 3.185 0.835 ;
        RECT  2.940 0.960 3.090 1.080 ;
        RECT  2.850 1.440 3.090 1.560 ;
        RECT  2.700 1.200 2.970 1.320 ;
        RECT  2.820 0.645 2.940 1.080 ;
        RECT  2.730 1.440 2.850 1.735 ;
        RECT  2.630 0.645 2.820 0.765 ;
        RECT  2.590 1.615 2.730 1.735 ;
        RECT  2.600 1.855 2.720 2.090 ;
        RECT  2.580 0.885 2.700 1.320 ;
        RECT  1.050 1.855 2.600 1.975 ;
        RECT  2.095 0.885 2.580 1.005 ;
        RECT  1.890 1.615 2.170 1.735 ;
        RECT  1.925 0.575 2.095 1.005 ;
        RECT  1.890 0.885 1.925 1.005 ;
        RECT  1.770 0.885 1.890 1.735 ;
        RECT  1.250 1.285 1.770 1.405 ;
        RECT  1.240 0.600 1.420 0.720 ;
        RECT  1.170 1.525 1.340 1.720 ;
        RECT  1.130 1.145 1.250 1.405 ;
        RECT  1.120 0.600 1.240 1.025 ;
        RECT  1.010 1.525 1.170 1.645 ;
        RECT  1.010 0.905 1.120 1.025 ;
        RECT  0.770 1.765 1.050 1.975 ;
        RECT  0.890 0.905 1.010 1.645 ;
        RECT  0.840 0.355 0.960 0.785 ;
        RECT  0.770 0.665 0.840 0.785 ;
        RECT  0.650 0.665 0.770 1.975 ;
        RECT  0.530 0.425 0.670 0.545 ;
        RECT  0.410 0.425 0.530 1.805 ;
    END
END MXI4XLAD
MACRO NAND2BX1AD
    CLASS CORE ;
    FOREIGN NAND2BX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.205 0.585 1.330 1.615 ;
        RECT  1.170 0.585 1.205 0.845 ;
        RECT  0.955 1.495 1.205 1.615 ;
        RECT  0.785 1.495 0.955 1.955 ;
        END
        AntennaDiffArea 0.23 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.865 0.780 1.375 ;
        END
        AntennaGateArea 0.091 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.865 0.490 1.225 ;
        END
        AntennaGateArea 0.042 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.635 -0.210 1.400 0.210 ;
        RECT  0.465 -0.210 0.635 0.505 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.315 2.310 1.400 2.730 ;
        RECT  1.145 1.785 1.315 2.730 ;
        RECT  0.565 2.310 1.145 2.730 ;
        RECT  0.395 1.825 0.565 2.730 ;
        RECT  0.000 2.310 0.395 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  1.020 1.020 1.085 1.280 ;
        RECT  0.900 0.625 1.020 1.280 ;
        RECT  0.255 0.625 0.900 0.745 ;
        RECT  0.190 0.575 0.255 0.745 ;
        RECT  0.190 1.375 0.255 1.545 ;
        RECT  0.070 0.575 0.190 1.545 ;
    END
END NAND2BX1AD
MACRO NAND2BX2AD
    CLASS CORE ;
    FOREIGN NAND2BX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.205 0.380 1.330 1.615 ;
        RECT  1.165 0.380 1.205 0.900 ;
        RECT  0.935 1.495 1.205 1.615 ;
        RECT  0.765 1.495 0.935 1.955 ;
        END
        AntennaDiffArea 0.435 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.865 0.775 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.865 0.490 1.225 ;
        END
        AntennaGateArea 0.0654 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.635 -0.210 1.400 0.210 ;
        RECT  0.465 -0.210 0.635 0.415 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.295 2.310 1.400 2.730 ;
        RECT  1.125 1.845 1.295 2.730 ;
        RECT  0.575 2.310 1.125 2.730 ;
        RECT  0.405 2.105 0.575 2.730 ;
        RECT  0.000 2.310 0.405 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  1.020 1.020 1.085 1.280 ;
        RECT  0.900 0.575 1.020 1.280 ;
        RECT  0.190 0.575 0.900 0.745 ;
        RECT  0.190 1.375 0.265 1.545 ;
        RECT  0.070 0.575 0.190 1.545 ;
    END
END NAND2BX2AD
MACRO NAND2BX4AD
    CLASS CORE ;
    FOREIGN NAND2BX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.795 2.170 1.655 ;
        RECT  1.345 0.795 2.010 0.925 ;
        RECT  1.705 1.525 2.010 1.655 ;
        RECT  1.535 1.525 1.705 2.055 ;
        RECT  0.985 1.525 1.535 1.655 ;
        RECT  1.175 0.410 1.345 0.925 ;
        RECT  0.815 1.525 0.985 2.060 ;
        END
        AntennaDiffArea 0.664 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.045 1.890 1.405 ;
        RECT  0.790 1.285 1.770 1.405 ;
        RECT  0.630 1.040 0.790 1.405 ;
        END
        AntennaGateArea 0.3249 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.055 0.270 1.225 ;
        RECT  0.070 1.055 0.210 1.485 ;
        END
        AntennaGateArea 0.129 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.005 -0.210 2.240 0.210 ;
        RECT  1.835 -0.210 2.005 0.675 ;
        RECT  0.680 -0.210 1.835 0.210 ;
        RECT  0.510 -0.210 0.680 0.675 ;
        RECT  0.000 -0.210 0.510 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.065 2.310 2.240 2.730 ;
        RECT  1.895 1.845 2.065 2.730 ;
        RECT  1.345 2.310 1.895 2.730 ;
        RECT  1.175 1.845 1.345 2.730 ;
        RECT  0.625 2.310 1.175 2.730 ;
        RECT  0.455 1.845 0.625 2.730 ;
        RECT  0.000 2.310 0.455 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.055 1.045 1.530 1.165 ;
        RECT  0.935 0.795 1.055 1.165 ;
        RECT  0.510 0.795 0.935 0.915 ;
        RECT  0.390 0.795 0.510 1.725 ;
        RECT  0.360 0.795 0.390 0.915 ;
        RECT  0.265 1.605 0.390 1.725 ;
        RECT  0.100 0.350 0.360 0.915 ;
        RECT  0.095 1.605 0.265 2.060 ;
    END
END NAND2BX4AD
MACRO NAND2BX8AD
    CLASS CORE ;
    FOREIGN NAND2BX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 0.480 3.820 1.795 ;
        RECT  3.110 0.480 3.610 0.730 ;
        RECT  3.450 1.330 3.610 1.795 ;
        RECT  3.245 1.330 3.450 2.075 ;
        RECT  3.230 1.555 3.245 2.075 ;
        RECT  2.730 1.555 3.230 1.795 ;
        RECT  2.850 0.350 3.110 0.730 ;
        RECT  1.670 0.480 2.850 0.730 ;
        RECT  2.510 1.555 2.730 2.100 ;
        RECT  2.015 1.555 2.510 1.795 ;
        RECT  1.795 1.555 2.015 2.100 ;
        RECT  1.285 1.555 1.795 1.795 ;
        RECT  1.410 0.350 1.670 0.730 ;
        RECT  1.075 1.555 1.285 2.100 ;
        END
        AntennaDiffArea 1.324 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.370 0.950 3.490 1.210 ;
        RECT  3.290 0.950 3.370 1.070 ;
        RECT  3.170 0.900 3.290 1.070 ;
        RECT  2.570 0.900 3.170 1.020 ;
        RECT  2.050 0.900 2.570 1.140 ;
        RECT  1.985 0.900 2.050 1.050 ;
        RECT  1.180 0.900 1.985 1.020 ;
        RECT  0.920 0.900 1.180 1.140 ;
        END
        AntennaGateArea 0.645 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.255 1.050 0.535 1.385 ;
        END
        AntennaGateArea 0.2597 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.795 -0.210 3.920 0.210 ;
        RECT  3.625 -0.210 3.795 0.360 ;
        RECT  2.335 -0.210 3.625 0.210 ;
        RECT  2.165 -0.210 2.335 0.360 ;
        RECT  1.015 -0.210 2.165 0.210 ;
        RECT  0.845 -0.210 1.015 0.675 ;
        RECT  0.265 -0.210 0.845 0.210 ;
        RECT  0.095 -0.210 0.265 0.675 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.785 2.310 3.920 2.730 ;
        RECT  3.615 1.975 3.785 2.730 ;
        RECT  3.065 2.310 3.615 2.730 ;
        RECT  2.895 1.975 3.065 2.730 ;
        RECT  2.345 2.310 2.895 2.730 ;
        RECT  2.175 1.975 2.345 2.730 ;
        RECT  1.625 2.310 2.175 2.730 ;
        RECT  1.455 1.975 1.625 2.730 ;
        RECT  0.905 2.310 1.455 2.730 ;
        RECT  0.735 1.825 0.905 2.730 ;
        RECT  0.255 2.310 0.735 2.730 ;
        RECT  0.085 2.205 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  2.770 1.140 3.030 1.385 ;
        RECT  1.635 1.265 2.770 1.385 ;
        RECT  1.375 1.140 1.635 1.385 ;
        RECT  0.800 1.265 1.375 1.385 ;
        RECT  0.680 0.795 0.800 1.635 ;
        RECT  0.670 0.795 0.680 0.915 ;
        RECT  0.545 1.515 0.680 1.635 ;
        RECT  0.550 0.350 0.670 0.915 ;
        RECT  0.410 0.350 0.550 0.730 ;
        RECT  0.375 1.515 0.545 1.945 ;
    END
END NAND2BX8AD
MACRO NAND2BXLAD
    CLASS CORE ;
    FOREIGN NAND2BXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.205 0.530 1.330 1.615 ;
        RECT  1.170 0.530 1.205 0.815 ;
        RECT  0.955 1.495 1.205 1.615 ;
        RECT  0.785 1.495 0.955 1.705 ;
        END
        AntennaDiffArea 0.15 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.625 0.865 0.780 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.865 0.490 1.225 ;
        END
        AntennaGateArea 0.0404 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.635 -0.210 1.400 0.210 ;
        RECT  0.465 -0.210 0.635 0.505 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.315 2.310 1.400 2.730 ;
        RECT  1.145 1.735 1.315 2.730 ;
        RECT  0.575 2.310 1.145 2.730 ;
        RECT  0.405 1.965 0.575 2.730 ;
        RECT  0.000 2.310 0.405 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  1.050 1.060 1.080 1.320 ;
        RECT  0.930 0.625 1.050 1.320 ;
        RECT  0.255 0.625 0.930 0.745 ;
        RECT  0.190 0.575 0.255 0.745 ;
        RECT  0.190 1.535 0.255 1.705 ;
        RECT  0.070 0.575 0.190 1.705 ;
    END
END NAND2BXLAD
MACRO NAND2X1AD
    CLASS CORE ;
    FOREIGN NAND2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 0.605 1.050 1.630 ;
        RECT  0.680 0.605 0.890 0.725 ;
        RECT  0.645 1.510 0.890 1.630 ;
        RECT  0.475 1.510 0.645 1.940 ;
        END
        AntennaDiffArea 0.233 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.035 0.405 1.205 ;
        RECT  0.070 1.035 0.210 1.655 ;
        END
        AntennaGateArea 0.09 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 0.845 0.770 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.285 -0.210 1.120 0.210 ;
        RECT  0.115 -0.210 0.285 0.830 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.005 2.310 1.120 2.730 ;
        RECT  0.835 1.750 1.005 2.730 ;
        RECT  0.285 2.310 0.835 2.730 ;
        RECT  0.115 1.775 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
	 END
END NAND2X1AD
MACRO NAND2X2AD
    CLASS CORE ;
    FOREIGN NAND2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 0.590 1.050 1.655 ;
        RECT  0.910 0.330 0.950 1.655 ;
        RECT  0.690 0.330 0.910 0.745 ;
        RECT  0.655 1.495 0.910 1.655 ;
        RECT  0.485 1.495 0.655 2.185 ;
        END
        AntennaDiffArea 0.401 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.010 0.240 1.655 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 0.865 0.770 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.295 -0.210 1.120 0.210 ;
        RECT  0.125 -0.210 0.295 0.755 ;
        RECT  0.000 -0.210 0.125 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.015 2.310 1.120 2.730 ;
        RECT  0.845 1.845 1.015 2.730 ;
        RECT  0.295 2.310 0.845 2.730 ;
        RECT  0.125 1.845 0.295 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
	 END
END NAND2X2AD
MACRO NAND2X3AD
    CLASS CORE ;
    FOREIGN NAND2X3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 0.835 1.890 1.675 ;
        RECT  1.065 0.835 1.730 0.955 ;
        RECT  1.425 1.555 1.730 1.675 ;
        RECT  1.255 1.555 1.425 2.060 ;
        RECT  0.705 1.555 1.255 1.675 ;
        RECT  0.895 0.345 1.065 0.955 ;
        RECT  0.535 1.555 0.705 2.060 ;
        END
        AntennaDiffArea 0.5 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.490 1.085 1.610 1.435 ;
        RECT  0.240 1.315 1.490 1.435 ;
        RECT  0.070 1.010 0.240 1.655 ;
        END
        AntennaGateArea 0.244 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.075 1.250 1.195 ;
        RECT  0.630 0.585 0.770 1.195 ;
        END
        AntennaGateArea 0.244 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.210 1.960 0.210 ;
        RECT  1.555 -0.210 1.725 0.715 ;
        RECT  0.405 -0.210 1.555 0.210 ;
        RECT  0.235 -0.210 0.405 0.715 ;
        RECT  0.000 -0.210 0.235 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.785 2.310 1.960 2.730 ;
        RECT  1.615 1.795 1.785 2.730 ;
        RECT  1.065 2.310 1.615 2.730 ;
        RECT  0.895 1.795 1.065 2.730 ;
        RECT  0.345 2.310 0.895 2.730 ;
        RECT  0.175 1.795 0.345 2.730 ;
        RECT  0.000 2.310 0.175 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
	 END
END NAND2X3AD
MACRO NAND2X4AD
    CLASS CORE ;
    FOREIGN NAND2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 0.795 1.890 1.655 ;
        RECT  1.065 0.795 1.730 0.925 ;
        RECT  1.425 1.525 1.730 1.655 ;
        RECT  1.255 1.525 1.425 2.055 ;
        RECT  0.705 1.525 1.255 1.655 ;
        RECT  0.895 0.410 1.065 0.925 ;
        RECT  0.535 1.525 0.705 2.060 ;
        END
        AntennaDiffArea 0.664 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 1.085 1.605 1.405 ;
        RECT  0.240 1.285 1.435 1.405 ;
        RECT  0.070 1.010 0.240 1.655 ;
        END
        AntennaGateArea 0.3249 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.045 1.250 1.165 ;
        RECT  0.630 0.585 0.770 1.165 ;
        END
        AntennaGateArea 0.324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.725 -0.210 1.960 0.210 ;
        RECT  1.555 -0.210 1.725 0.675 ;
        RECT  0.405 -0.210 1.555 0.210 ;
        RECT  0.235 -0.210 0.405 0.790 ;
        RECT  0.000 -0.210 0.235 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.785 2.310 1.960 2.730 ;
        RECT  1.615 1.775 1.785 2.730 ;
        RECT  1.065 2.310 1.615 2.730 ;
        RECT  0.895 1.775 1.065 2.730 ;
        RECT  0.345 2.310 0.895 2.730 ;
        RECT  0.175 1.775 0.345 2.730 ;
        RECT  0.000 2.310 0.175 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
	 END
END NAND2X4AD
MACRO NAND2X5AD
    CLASS CORE ;
    FOREIGN NAND2X5AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.375 0.570 2.450 1.695 ;
        RECT  2.280 0.355 2.375 1.695 ;
        RECT  2.205 0.355 2.280 0.785 ;
        RECT  2.075 1.545 2.280 1.695 ;
        RECT  0.995 0.570 2.205 0.745 ;
        RECT  1.905 1.545 2.075 2.010 ;
        RECT  1.355 1.545 1.905 1.695 ;
        RECT  1.185 1.545 1.355 2.010 ;
        RECT  0.635 1.545 1.185 1.695 ;
        RECT  0.825 0.340 0.995 0.770 ;
        RECT  0.465 1.545 0.635 2.035 ;
        END
        AntennaDiffArea 0.889 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 0.985 1.620 1.105 ;
        RECT  1.260 0.890 1.380 1.105 ;
        RECT  0.235 0.890 1.260 1.010 ;
        RECT  0.070 0.890 0.235 1.655 ;
        END
        AntennaGateArea 0.408 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.005 2.150 1.265 ;
        RECT  1.750 0.865 1.890 1.375 ;
        RECT  1.000 1.255 1.750 1.375 ;
        RECT  0.830 1.130 1.000 1.375 ;
        END
        AntennaGateArea 0.408 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.665 -0.210 2.520 0.210 ;
        RECT  1.495 -0.210 1.665 0.415 ;
        RECT  0.335 -0.210 1.495 0.210 ;
        RECT  0.165 -0.210 0.335 0.675 ;
        RECT  0.000 -0.210 0.165 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 2.310 2.520 2.730 ;
        RECT  2.265 1.845 2.435 2.730 ;
        RECT  1.715 2.310 2.265 2.730 ;
        RECT  1.545 1.845 1.715 2.730 ;
        RECT  0.995 2.310 1.545 2.730 ;
        RECT  0.825 1.845 0.995 2.730 ;
        RECT  0.275 2.310 0.825 2.730 ;
        RECT  0.105 1.845 0.275 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
	 END
END NAND2X5AD
MACRO NAND2X6AD
    CLASS CORE ;
    FOREIGN NAND2X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.325 0.570 2.450 1.725 ;
        RECT  2.285 0.340 2.325 1.725 ;
        RECT  2.155 0.340 2.285 0.770 ;
        RECT  2.075 1.550 2.285 1.725 ;
        RECT  0.995 0.570 2.155 0.745 ;
        RECT  1.905 1.550 2.075 2.010 ;
        RECT  1.355 1.550 1.905 1.725 ;
        RECT  1.185 1.550 1.355 2.010 ;
        RECT  0.635 1.550 1.185 1.725 ;
        RECT  0.825 0.340 0.995 0.770 ;
        RECT  0.465 1.550 0.635 2.015 ;
        END
        AntennaDiffArea 1.065 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.020 1.620 1.140 ;
        RECT  1.260 0.890 1.380 1.140 ;
        RECT  0.235 0.890 1.260 1.010 ;
        RECT  0.070 0.890 0.235 1.655 ;
        END
        AntennaGateArea 0.486 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.005 2.150 1.265 ;
        RECT  1.750 0.865 1.890 1.380 ;
        RECT  1.045 1.260 1.750 1.380 ;
        RECT  0.785 1.130 1.045 1.380 ;
        END
        AntennaGateArea 0.486 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.665 -0.210 2.520 0.210 ;
        RECT  1.495 -0.210 1.665 0.415 ;
        RECT  0.385 -0.210 1.495 0.210 ;
        RECT  0.215 -0.210 0.385 0.675 ;
        RECT  0.000 -0.210 0.215 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.435 2.310 2.520 2.730 ;
        RECT  2.265 1.845 2.435 2.730 ;
        RECT  1.715 2.310 2.265 2.730 ;
        RECT  1.545 1.845 1.715 2.730 ;
        RECT  0.995 2.310 1.545 2.730 ;
        RECT  0.825 1.845 0.995 2.730 ;
        RECT  0.275 2.310 0.825 2.730 ;
        RECT  0.105 1.845 0.275 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
	 END
END NAND2X6AD
MACRO NAND2X8AD
    CLASS CORE ;
    FOREIGN NAND2X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 0.480 3.260 2.075 ;
        RECT  2.460 0.480 3.010 0.730 ;
        RECT  2.615 1.555 3.010 2.075 ;
        RECT  2.090 1.555 2.615 1.795 ;
        RECT  2.200 0.350 2.460 0.730 ;
        RECT  1.030 0.480 2.200 0.730 ;
        RECT  1.870 1.555 2.090 2.100 ;
        RECT  1.375 1.555 1.870 1.795 ;
        RECT  1.155 1.555 1.375 2.100 ;
        RECT  0.645 1.555 1.155 1.795 ;
        RECT  0.770 0.350 1.030 0.730 ;
        RECT  0.435 1.555 0.645 2.100 ;
        END
        AntennaDiffArea 1.328 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.730 0.990 2.850 1.250 ;
        RECT  2.610 0.900 2.730 1.110 ;
        RECT  1.945 0.900 2.610 1.020 ;
        RECT  1.425 0.900 1.945 1.140 ;
        RECT  0.405 0.900 1.425 1.020 ;
        RECT  0.235 0.900 0.405 1.195 ;
        END
        AntennaGateArea 0.648 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 1.140 2.470 1.385 ;
        RECT  1.095 1.265 2.210 1.385 ;
        RECT  0.585 1.140 1.095 1.385 ;
        END
        AntennaGateArea 0.6489 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.095 -0.210 3.360 0.210 ;
        RECT  2.925 -0.210 3.095 0.360 ;
        RECT  1.700 -0.210 2.925 0.210 ;
        RECT  1.530 -0.210 1.700 0.360 ;
        RECT  0.375 -0.210 1.530 0.210 ;
        RECT  0.205 -0.210 0.375 0.675 ;
        RECT  0.000 -0.210 0.205 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.215 2.310 3.360 2.730 ;
        RECT  3.045 2.195 3.215 2.730 ;
        RECT  2.425 2.310 3.045 2.730 ;
        RECT  2.255 1.975 2.425 2.730 ;
        RECT  1.705 2.310 2.255 2.730 ;
        RECT  1.535 1.975 1.705 2.730 ;
        RECT  0.985 2.310 1.535 2.730 ;
        RECT  0.815 1.975 0.985 2.730 ;
        RECT  0.265 2.310 0.815 2.730 ;
        RECT  0.095 1.530 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
	 END
END NAND2X8AD
MACRO NAND2XLAD
    CLASS CORE ;
    FOREIGN NAND2XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.600 1.050 1.615 ;
        RECT  0.720 0.600 0.910 0.720 ;
        RECT  0.625 1.495 0.910 1.615 ;
        RECT  0.455 1.495 0.625 1.785 ;
        END
        AntennaDiffArea 0.161 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.165 0.865 0.335 1.350 ;
        RECT  0.070 0.865 0.165 1.095 ;
        END
        AntennaGateArea 0.06 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.605 0.865 0.790 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.255 -0.210 1.120 0.210 ;
        RECT  0.085 -0.210 0.255 0.745 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.985 2.310 1.120 2.730 ;
        RECT  0.815 1.735 0.985 2.730 ;
        RECT  0.265 2.310 0.815 2.730 ;
        RECT  0.095 1.735 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
	 END
END NAND2XLAD
MACRO NAND3BX1AD
    CLASS CORE ;
    FOREIGN NAND3BX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.595 0.450 1.610 1.630 ;
        RECT  1.470 0.450 1.595 1.940 ;
        RECT  1.425 0.450 1.470 0.620 ;
        RECT  1.425 1.510 1.470 1.940 ;
        RECT  0.925 1.510 1.425 1.630 ;
        RECT  0.755 1.510 0.925 1.940 ;
        END
        AntennaDiffArea 0.365 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.770 1.375 ;
        END
        AntennaGateArea 0.0904 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.0904 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.500 1.375 ;
        RECT  0.325 0.865 0.350 1.125 ;
        END
        AntennaGateArea 0.0414 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.670 -0.210 1.680 0.210 ;
        RECT  0.410 -0.210 0.670 0.505 ;
        RECT  0.000 -0.210 0.410 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.180 2.310 1.680 2.730 ;
        RECT  0.490 2.215 1.180 2.730 ;
        RECT  0.000 2.310 0.490 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.290 0.960 1.350 1.220 ;
        RECT  1.170 0.625 1.290 1.220 ;
        RECT  0.255 0.625 1.170 0.745 ;
        RECT  0.205 0.360 0.255 0.745 ;
        RECT  0.205 1.340 0.230 1.600 ;
        RECT  0.085 0.360 0.205 1.600 ;
    END
END NAND3BX1AD
MACRO NAND3BX2AD
    CLASS CORE ;
    FOREIGN NAND3BX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.805 0.665 1.890 1.725 ;
        RECT  1.750 0.665 1.805 2.030 ;
        RECT  1.735 0.665 1.750 0.805 ;
        RECT  1.635 1.585 1.750 2.030 ;
        RECT  1.565 0.360 1.735 0.805 ;
        RECT  1.085 1.585 1.635 1.725 ;
        RECT  0.915 1.585 1.085 2.030 ;
        END
        AntennaDiffArea 0.615 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.845 1.215 ;
        END
        AntennaGateArea 0.162 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.080 0.585 1.330 1.215 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.045 0.270 1.215 ;
        RECT  0.070 1.045 0.210 1.435 ;
        END
        AntennaGateArea 0.0654 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.725 -0.210 1.960 0.210 ;
        RECT  0.555 -0.210 0.725 0.675 ;
        RECT  0.000 -0.210 0.555 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.445 2.310 1.960 2.730 ;
        RECT  1.275 1.845 1.445 2.730 ;
        RECT  0.725 2.310 1.275 2.730 ;
        RECT  0.555 1.840 0.725 2.730 ;
        RECT  0.000 2.310 0.555 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.450 1.020 1.570 1.465 ;
        RECT  0.510 1.345 1.450 1.465 ;
        RECT  0.390 0.795 0.510 1.675 ;
        RECT  0.345 0.795 0.390 0.915 ;
        RECT  0.345 1.555 0.390 1.675 ;
        RECT  0.175 0.665 0.345 0.915 ;
        RECT  0.175 1.555 0.345 1.725 ;
    END
END NAND3BX2AD
MACRO NAND3BX4AD
    CLASS CORE ;
    FOREIGN NAND3BX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.430 0.630 2.590 1.720 ;
        RECT  1.880 0.630 2.430 0.805 ;
        RECT  0.905 1.550 2.430 1.720 ;
        RECT  1.710 0.375 1.880 0.805 ;
        END
        AntennaDiffArea 0.962 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.710 1.000 2.830 2.010 ;
        RECT  0.770 1.890 2.710 2.010 ;
        RECT  0.630 1.020 0.770 2.010 ;
        END
        AntennaGateArea 0.324 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 1.010 2.310 1.400 ;
        RECT  1.330 1.280 2.190 1.400 ;
        RECT  1.190 0.865 1.330 1.400 ;
        END
        AntennaGateArea 0.324 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.240 1.375 ;
        END
        AntennaGateArea 0.1294 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.870 -0.210 3.080 0.210 ;
        RECT  2.710 -0.210 2.870 0.875 ;
        RECT  0.850 -0.210 2.710 0.210 ;
        RECT  0.590 -0.210 0.850 0.505 ;
        RECT  0.000 -0.210 0.590 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.980 2.310 3.080 2.730 ;
        RECT  2.720 2.130 2.980 2.730 ;
        RECT  2.260 2.310 2.720 2.730 ;
        RECT  2.000 2.130 2.260 2.730 ;
        RECT  1.540 2.310 2.000 2.730 ;
        RECT  1.280 2.130 1.540 2.730 ;
        RECT  0.740 2.310 1.280 2.730 ;
        RECT  0.480 2.130 0.740 2.730 ;
        RECT  0.000 2.310 0.480 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  1.570 1.040 2.045 1.160 ;
        RECT  1.450 0.625 1.570 1.160 ;
        RECT  0.490 0.625 1.450 0.745 ;
        RECT  0.370 0.625 0.490 1.680 ;
        RECT  0.345 0.625 0.370 0.745 ;
        RECT  0.315 1.560 0.370 1.680 ;
        RECT  0.175 0.560 0.345 0.745 ;
        RECT  0.145 1.560 0.315 1.990 ;
    END
END NAND3BX4AD
MACRO NAND3BXLAD
    CLASS CORE ;
    FOREIGN NAND3BXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.360 1.610 1.680 ;
        RECT  1.425 0.360 1.470 0.530 ;
        RECT  1.425 1.510 1.470 1.680 ;
        RECT  0.925 1.510 1.425 1.630 ;
        RECT  0.755 1.510 0.925 1.680 ;
        END
        AntennaDiffArea 0.242 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.770 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.500 1.375 ;
        RECT  0.325 0.865 0.350 1.125 ;
        END
        AntennaGateArea 0.0404 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.670 -0.210 1.680 0.210 ;
        RECT  0.410 -0.210 0.670 0.505 ;
        RECT  0.000 -0.210 0.410 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.215 2.310 1.680 2.730 ;
        RECT  1.045 2.005 1.215 2.730 ;
        RECT  0.635 2.310 1.045 2.730 ;
        RECT  0.465 2.005 0.635 2.730 ;
        RECT  0.000 2.310 0.465 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.290 0.960 1.350 1.220 ;
        RECT  1.170 0.625 1.290 1.220 ;
        RECT  0.255 0.625 1.170 0.745 ;
        RECT  0.205 0.360 0.255 0.745 ;
        RECT  0.205 1.330 0.230 1.590 ;
        RECT  0.085 0.360 0.205 1.590 ;
    END
END NAND3BXLAD
MACRO NAND3X1AD
    CLASS CORE ;
    FOREIGN NAND3X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.315 0.605 1.330 1.630 ;
        RECT  1.190 0.605 1.315 1.940 ;
        RECT  1.000 0.605 1.190 0.725 ;
        RECT  1.145 1.510 1.190 1.940 ;
        RECT  0.595 1.510 1.145 1.630 ;
        RECT  0.425 1.510 0.595 1.940 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.035 0.425 1.205 ;
        RECT  0.070 1.035 0.210 1.655 ;
        END
        AntennaGateArea 0.0904 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 0.845 0.770 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.255 -0.210 1.400 0.210 ;
        RECT  0.085 -0.210 0.255 0.750 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.955 2.310 1.400 2.730 ;
        RECT  0.785 1.750 0.955 2.730 ;
        RECT  0.255 2.310 0.785 2.730 ;
        RECT  0.085 2.215 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
	 END
END NAND3X1AD
MACRO NAND3X2AD
    CLASS CORE ;
    FOREIGN NAND3X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.265 1.510 1.435 1.955 ;
        RECT  1.145 0.430 1.315 0.875 ;
        RECT  1.050 1.510 1.265 1.650 ;
        RECT  1.050 0.705 1.145 0.875 ;
        RECT  0.910 0.705 1.050 1.650 ;
        RECT  0.715 1.510 0.910 1.650 ;
        RECT  0.545 1.510 0.715 1.955 ;
        END
        AntennaDiffArea 0.615 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.000 0.480 1.375 ;
        RECT  0.070 1.145 0.320 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.780 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.140 1.610 1.375 ;
        RECT  1.190 1.020 1.350 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.360 -0.210 1.680 0.210 ;
        RECT  0.180 -0.210 0.360 0.675 ;
        RECT  0.000 -0.210 0.180 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.075 2.310 1.680 2.730 ;
        RECT  0.905 1.775 1.075 2.730 ;
        RECT  0.355 2.310 0.905 2.730 ;
        RECT  0.185 1.515 0.355 2.730 ;
        RECT  0.000 2.310 0.185 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
	 END
END NAND3X2AD
MACRO NAND3X3AD
    CLASS CORE ;
    FOREIGN NAND3X3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.515 2.100 1.635 ;
        RECT  1.050 0.620 1.275 0.790 ;
        RECT  0.910 0.620 1.050 1.635 ;
        RECT  0.400 1.515 0.910 1.635 ;
        END
        AntennaDiffArea 0.718 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.225 1.195 2.345 1.875 ;
        RECT  2.150 1.195 2.225 1.315 ;
        RECT  0.230 1.755 2.225 1.875 ;
        RECT  2.030 1.000 2.150 1.315 ;
        RECT  0.070 0.865 0.230 1.875 ;
        END
        AntennaGateArea 0.246 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 0.380 1.850 1.265 ;
        RECT  0.770 0.380 1.730 0.500 ;
        RECT  0.620 0.380 0.770 1.375 ;
        END
        AntennaGateArea 0.246 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.145 1.610 1.375 ;
        RECT  1.170 0.910 1.330 1.375 ;
        END
        AntennaGateArea 0.246 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.210 2.520 0.210 ;
        RECT  2.150 -0.210 2.330 0.730 ;
        RECT  0.320 -0.210 2.150 0.210 ;
        RECT  0.140 -0.210 0.320 0.730 ;
        RECT  0.000 -0.210 0.140 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.415 2.310 2.520 2.730 ;
        RECT  2.245 1.995 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 1.995 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.995 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.995 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
	 END
END NAND3X3AD
MACRO NAND3X4AD
    CLASS CORE ;
    FOREIGN NAND3X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.495 2.055 1.665 ;
        RECT  1.050 0.620 1.275 0.790 ;
        RECT  0.910 0.620 1.050 1.665 ;
        RECT  0.445 1.495 0.910 1.665 ;
        END
        AntennaDiffArea 0.946 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.215 1.195 2.335 1.955 ;
        RECT  2.150 1.195 2.215 1.315 ;
        RECT  0.230 1.835 2.215 1.955 ;
        RECT  2.030 1.000 2.150 1.315 ;
        RECT  0.070 0.865 0.230 1.955 ;
        END
        AntennaGateArea 0.324 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 0.380 1.850 1.265 ;
        RECT  0.770 0.380 1.730 0.500 ;
        RECT  0.620 0.380 0.770 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.145 1.610 1.375 ;
        RECT  1.170 0.910 1.330 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.330 -0.210 2.520 0.210 ;
        RECT  2.150 -0.210 2.330 0.675 ;
        RECT  0.320 -0.210 2.150 0.210 ;
        RECT  0.140 -0.210 0.320 0.675 ;
        RECT  0.000 -0.210 0.140 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.415 2.310 2.520 2.730 ;
        RECT  2.245 2.075 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 2.075 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 2.075 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 2.075 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
	 END
END NAND3X4AD
MACRO NAND3X6AD
    CLASS CORE ;
    FOREIGN NAND3X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.540 0.585 3.570 1.375 ;
        RECT  3.445 0.585 3.540 1.985 ;
        RECT  3.400 0.330 3.445 1.985 ;
        RECT  3.275 0.330 3.400 0.760 ;
        RECT  3.325 1.375 3.400 1.985 ;
        RECT  0.615 1.815 3.325 1.985 ;
        RECT  2.260 0.455 3.275 0.635 ;
        RECT  2.120 0.380 2.260 0.635 ;
        RECT  1.060 0.380 2.120 0.520 ;
        RECT  0.445 1.540 0.615 1.985 ;
        END
        AntennaDiffArea 1.561 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.040 2.510 1.160 ;
        RECT  1.880 0.640 2.000 1.160 ;
        RECT  0.230 0.640 1.880 0.760 ;
        RECT  0.070 0.640 0.230 1.375 ;
        END
        AntennaGateArea 0.486 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.780 1.005 2.900 1.400 ;
        RECT  1.760 1.280 2.780 1.400 ;
        RECT  1.640 0.880 1.760 1.400 ;
        RECT  0.770 0.880 1.640 1.000 ;
        RECT  0.620 0.880 0.770 1.375 ;
        END
        AntennaGateArea 0.486 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.080 1.005 3.200 1.670 ;
        RECT  1.330 1.550 3.080 1.670 ;
        RECT  1.330 1.120 1.460 1.240 ;
        RECT  1.190 1.120 1.330 1.670 ;
        RECT  0.940 1.120 1.190 1.240 ;
        END
        AntennaGateArea 0.486 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.395 -0.210 3.640 0.210 ;
        RECT  2.225 -0.210 2.395 0.260 ;
        RECT  0.320 -0.210 2.225 0.210 ;
        RECT  0.140 -0.210 0.320 0.415 ;
        RECT  0.000 -0.210 0.140 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.135 2.310 3.640 2.730 ;
        RECT  2.965 2.105 3.135 2.730 ;
        RECT  2.415 2.310 2.965 2.730 ;
        RECT  2.245 2.105 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 2.105 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 2.105 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.585 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
	 END
END NAND3X6AD
MACRO NAND3X8AD
    CLASS CORE ;
    FOREIGN NAND3X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.460 0.380 4.660 2.075 ;
        RECT  1.060 0.380 4.460 0.520 ;
        RECT  4.130 1.505 4.460 2.075 ;
        RECT  4.045 1.505 4.130 2.010 ;
        RECT  3.495 1.810 4.045 2.010 ;
        RECT  3.325 1.505 3.495 2.010 ;
        RECT  0.615 1.810 3.325 2.010 ;
        RECT  0.445 1.540 0.615 2.010 ;
        END
        AntennaDiffArea 1.886 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.160 0.640 4.280 1.265 ;
        RECT  2.610 0.640 4.160 0.760 ;
        RECT  2.490 0.640 2.610 1.160 ;
        RECT  2.110 1.040 2.490 1.160 ;
        RECT  1.990 0.640 2.110 1.160 ;
        RECT  0.230 0.640 1.990 0.760 ;
        RECT  0.070 0.640 0.230 1.375 ;
        END
        AntennaGateArea 0.648 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.860 0.880 3.980 1.265 ;
        RECT  2.900 0.880 3.860 1.000 ;
        RECT  2.780 0.880 2.900 1.400 ;
        RECT  1.760 1.280 2.780 1.400 ;
        RECT  1.640 0.880 1.760 1.400 ;
        RECT  0.770 0.880 1.640 1.000 ;
        RECT  0.620 0.880 0.770 1.375 ;
        END
        AntennaGateArea 0.648 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.185 1.120 3.640 1.240 ;
        RECT  3.065 1.120 3.185 1.640 ;
        RECT  1.330 1.520 3.065 1.640 ;
        RECT  1.330 1.120 1.460 1.240 ;
        RECT  1.190 1.120 1.330 1.640 ;
        RECT  0.940 1.120 1.190 1.240 ;
        END
        AntennaGateArea 0.648 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.595 -0.210 4.760 0.210 ;
        RECT  4.425 -0.210 4.595 0.260 ;
        RECT  2.395 -0.210 4.425 0.210 ;
        RECT  2.225 -0.210 2.395 0.260 ;
        RECT  0.320 -0.210 2.225 0.210 ;
        RECT  0.140 -0.210 0.320 0.415 ;
        RECT  0.000 -0.210 0.140 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.645 2.310 4.760 2.730 ;
        RECT  4.475 2.195 4.645 2.730 ;
        RECT  3.900 2.310 4.475 2.730 ;
        RECT  3.640 2.130 3.900 2.730 ;
        RECT  3.180 2.310 3.640 2.730 ;
        RECT  2.920 2.130 3.180 2.730 ;
        RECT  2.460 2.310 2.920 2.730 ;
        RECT  2.200 2.130 2.460 2.730 ;
        RECT  1.740 2.310 2.200 2.730 ;
        RECT  1.480 2.130 1.740 2.730 ;
        RECT  1.020 2.310 1.480 2.730 ;
        RECT  0.760 2.130 1.020 2.730 ;
        RECT  0.255 2.310 0.760 2.730 ;
        RECT  0.085 1.585 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.760 2.520 ;
	 END
END NAND3X8AD
MACRO NAND3XLAD
    CLASS CORE ;
    FOREIGN NAND3XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.605 1.330 1.720 ;
        RECT  1.040 0.605 1.190 0.725 ;
        RECT  1.145 1.510 1.190 1.720 ;
        RECT  0.595 1.510 1.145 1.630 ;
        RECT  0.425 1.510 0.595 1.720 ;
        END
        AntennaDiffArea 0.246 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.035 0.415 1.205 ;
        RECT  0.070 1.035 0.210 1.655 ;
        END
        AntennaGateArea 0.0604 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 0.845 0.770 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.295 -0.210 1.400 0.210 ;
        RECT  0.125 -0.210 0.295 0.750 ;
        RECT  0.000 -0.210 0.125 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.955 2.310 1.400 2.730 ;
        RECT  0.785 1.750 0.955 2.730 ;
        RECT  0.255 2.310 0.785 2.730 ;
        RECT  0.085 2.180 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
	 END
END NAND3XLAD
MACRO NAND4BBX1AD
    CLASS CORE ;
    FOREIGN NAND4BBX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 0.645 2.730 1.615 ;
        RECT  2.355 1.495 2.570 1.615 ;
        RECT  2.185 1.495 2.355 2.015 ;
        RECT  1.635 1.495 2.185 1.615 ;
        RECT  1.465 1.495 1.635 2.015 ;
        END
        AntennaDiffArea 0.391 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.000 1.590 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.720 0.930 1.890 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.780 1.275 ;
        END
        AntennaGateArea 0.0414 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.010 0.235 1.375 ;
        END
        AntennaGateArea 0.0414 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.420 -0.210 2.800 0.210 ;
        RECT  1.160 -0.210 1.420 0.310 ;
        RECT  0.680 -0.210 1.160 0.210 ;
        RECT  0.420 -0.210 0.680 0.310 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.715 2.310 2.800 2.730 ;
        RECT  2.545 1.735 2.715 2.730 ;
        RECT  1.995 2.310 2.545 2.730 ;
        RECT  1.825 1.735 1.995 2.730 ;
        RECT  1.275 2.310 1.825 2.730 ;
        RECT  1.105 1.950 1.275 2.730 ;
        RECT  0.605 2.310 1.105 2.730 ;
        RECT  0.435 1.925 0.605 2.730 ;
        RECT  0.000 2.310 0.435 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.410 1.000 2.450 1.260 ;
        RECT  2.290 0.430 2.410 1.260 ;
        RECT  0.510 0.430 2.290 0.550 ;
        RECT  2.030 0.670 2.150 1.260 ;
        RECT  1.020 0.670 2.030 0.790 ;
        RECT  0.900 0.670 1.020 1.710 ;
        RECT  0.810 1.450 0.900 1.710 ;
        RECT  0.390 0.430 0.510 1.615 ;
        RECT  0.085 0.720 0.390 0.890 ;
        RECT  0.255 1.495 0.390 1.615 ;
        RECT  0.085 1.495 0.255 1.665 ;
    END
END NAND4BBX1AD
MACRO NAND4BBX2AD
    CLASS CORE ;
    FOREIGN NAND4BBX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 0.355 2.730 1.615 ;
        RECT  2.355 1.495 2.570 1.615 ;
        RECT  2.185 1.495 2.355 1.940 ;
        RECT  1.635 1.495 2.185 1.615 ;
        RECT  1.465 1.495 1.635 1.940 ;
        END
        AntennaDiffArea 0.663 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.000 1.590 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.720 0.930 1.890 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.780 1.275 ;
        END
        AntennaGateArea 0.0654 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.980 0.235 1.375 ;
        END
        AntennaGateArea 0.0654 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.370 -0.210 2.800 0.210 ;
        RECT  1.110 -0.210 1.370 0.310 ;
        RECT  0.680 -0.210 1.110 0.210 ;
        RECT  0.420 -0.210 0.680 0.310 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.715 2.310 2.800 2.730 ;
        RECT  2.545 1.845 2.715 2.730 ;
        RECT  1.995 2.310 2.545 2.730 ;
        RECT  1.825 1.845 1.995 2.730 ;
        RECT  1.275 2.310 1.825 2.730 ;
        RECT  1.105 1.950 1.275 2.730 ;
        RECT  0.605 2.310 1.105 2.730 ;
        RECT  0.435 1.985 0.605 2.730 ;
        RECT  0.000 2.310 0.435 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.410 1.000 2.450 1.260 ;
        RECT  2.290 0.430 2.410 1.260 ;
        RECT  0.510 0.430 2.290 0.550 ;
        RECT  2.030 0.670 2.150 1.260 ;
        RECT  1.020 0.670 2.030 0.790 ;
        RECT  0.900 0.670 1.020 1.710 ;
        RECT  0.810 1.450 0.900 1.710 ;
        RECT  0.390 0.430 0.510 1.615 ;
        RECT  0.085 0.685 0.390 0.855 ;
        RECT  0.255 1.495 0.390 1.615 ;
        RECT  0.085 1.495 0.255 1.665 ;
    END
END NAND4BBX2AD
MACRO NAND4BBX4AD
    CLASS CORE ;
    FOREIGN NAND4BBX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.270 0.710 4.410 1.570 ;
        RECT  2.865 0.710 4.270 0.840 ;
        RECT  4.130 1.440 4.270 1.570 ;
        RECT  4.010 1.440 4.130 2.130 ;
        RECT  1.490 2.000 4.010 2.130 ;
        RECT  2.695 0.410 2.865 0.840 ;
        END
        AntennaDiffArea 1.124 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.020 4.130 1.295 ;
        RECT  3.890 1.175 4.010 1.295 ;
        RECT  3.770 1.175 3.890 1.880 ;
        RECT  1.610 1.760 3.770 1.880 ;
        RECT  1.470 1.020 1.610 1.880 ;
        END
        AntennaGateArea 0.32 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.530 1.020 3.650 1.640 ;
        RECT  1.910 1.520 3.530 1.640 ;
        RECT  1.740 1.025 1.910 1.640 ;
        END
        AntennaGateArea 0.3224 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 0.865 0.770 1.375 ;
        END
        AntennaGateArea 0.129 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.240 1.260 ;
        END
        AntennaGateArea 0.129 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.305 -0.210 4.480 0.210 ;
        RECT  4.135 -0.210 4.305 0.535 ;
        RECT  1.440 -0.210 4.135 0.210 ;
        RECT  1.180 -0.210 1.440 0.330 ;
        RECT  0.690 -0.210 1.180 0.210 ;
        RECT  0.430 -0.210 0.690 0.330 ;
        RECT  0.000 -0.210 0.430 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.370 2.310 4.480 2.730 ;
        RECT  4.250 1.730 4.370 2.730 ;
        RECT  3.665 2.310 4.250 2.730 ;
        RECT  3.405 2.250 3.665 2.730 ;
        RECT  2.890 2.310 3.405 2.730 ;
        RECT  2.630 2.250 2.890 2.730 ;
        RECT  2.130 2.310 2.630 2.730 ;
        RECT  1.870 2.250 2.130 2.730 ;
        RECT  1.320 2.310 1.870 2.730 ;
        RECT  1.200 1.690 1.320 2.730 ;
        RECT  0.615 2.310 1.200 2.730 ;
        RECT  0.445 1.665 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
        LAYER M1 ;
        RECT  3.200 1.020 3.320 1.400 ;
        RECT  2.290 1.280 3.200 1.400 ;
        RECT  2.560 1.040 3.010 1.160 ;
        RECT  2.440 0.450 2.560 1.160 ;
        RECT  0.480 0.450 2.440 0.570 ;
        RECT  2.170 0.690 2.290 1.400 ;
        RECT  1.010 0.690 2.170 0.810 ;
        RECT  0.975 0.690 1.010 1.615 ;
        RECT  0.890 0.690 0.975 2.095 ;
        RECT  0.855 1.495 0.890 2.095 ;
        RECT  0.805 1.665 0.855 2.095 ;
        RECT  0.360 0.450 0.480 1.540 ;
        RECT  0.110 0.450 0.360 0.710 ;
        RECT  0.230 1.420 0.360 1.540 ;
        RECT  0.110 1.420 0.230 1.940 ;
    END
END NAND4BBX4AD
MACRO NAND4BBXLAD
    CLASS CORE ;
    FOREIGN NAND4BBXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 0.645 2.730 1.715 ;
        RECT  2.355 1.595 2.570 1.715 ;
        RECT  2.185 1.595 2.355 1.805 ;
        RECT  1.635 1.595 2.185 1.715 ;
        RECT  1.465 1.595 1.635 1.805 ;
        END
        AntennaDiffArea 0.26 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.000 1.590 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.720 0.930 1.890 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.780 1.275 ;
        END
        AntennaGateArea 0.0404 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.010 0.235 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.420 -0.210 2.800 0.210 ;
        RECT  1.160 -0.210 1.420 0.310 ;
        RECT  0.680 -0.210 1.160 0.210 ;
        RECT  0.420 -0.210 0.680 0.310 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.715 2.310 2.800 2.730 ;
        RECT  2.545 1.835 2.715 2.730 ;
        RECT  1.995 2.310 2.545 2.730 ;
        RECT  1.825 1.835 1.995 2.730 ;
        RECT  1.275 2.310 1.825 2.730 ;
        RECT  1.105 1.835 1.275 2.730 ;
        RECT  0.605 2.310 1.105 2.730 ;
        RECT  0.435 1.925 0.605 2.730 ;
        RECT  0.000 2.310 0.435 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.410 1.000 2.450 1.260 ;
        RECT  2.290 0.430 2.410 1.260 ;
        RECT  0.510 0.430 2.290 0.550 ;
        RECT  2.030 0.670 2.150 1.260 ;
        RECT  1.020 0.670 2.030 0.790 ;
        RECT  0.900 0.670 1.020 1.710 ;
        RECT  0.810 1.450 0.900 1.710 ;
        RECT  0.390 0.430 0.510 1.615 ;
        RECT  0.085 0.720 0.390 0.890 ;
        RECT  0.255 1.495 0.390 1.615 ;
        RECT  0.085 1.495 0.255 1.665 ;
    END
END NAND4BBXLAD
MACRO NAND4BX1AD
    CLASS CORE ;
    FOREIGN NAND4BX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.475 2.170 1.645 ;
        RECT  1.915 0.475 2.030 0.645 ;
        RECT  1.795 1.525 2.030 1.645 ;
        RECT  1.625 1.525 1.795 1.955 ;
        RECT  1.075 1.525 1.625 1.645 ;
        RECT  0.905 1.525 1.075 1.955 ;
        END
        AntennaDiffArea 0.391 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.770 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.995 1.200 1.255 ;
        RECT  0.910 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.410 1.005 1.610 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.235 1.375 ;
        END
        AntennaGateArea 0.0425 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.725 -0.210 2.240 0.210 ;
        RECT  0.555 -0.210 0.725 0.505 ;
        RECT  0.000 -0.210 0.555 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.155 2.310 2.240 2.730 ;
        RECT  1.985 1.815 2.155 2.730 ;
        RECT  1.435 2.310 1.985 2.730 ;
        RECT  1.265 1.815 1.435 2.730 ;
        RECT  0.715 2.310 1.265 2.730 ;
        RECT  0.545 1.815 0.715 2.730 ;
        RECT  0.000 2.310 0.545 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.790 0.765 1.910 1.130 ;
        RECT  1.720 0.765 1.790 0.885 ;
        RECT  1.600 0.625 1.720 0.885 ;
        RECT  0.510 0.625 1.600 0.745 ;
        RECT  0.390 0.625 0.510 1.625 ;
        RECT  0.335 0.625 0.390 0.745 ;
        RECT  0.335 1.505 0.390 1.625 ;
        RECT  0.165 0.565 0.335 0.745 ;
        RECT  0.165 1.505 0.335 1.675 ;
    END
END NAND4BX1AD
MACRO NAND4BX2AD
    CLASS CORE ;
    FOREIGN NAND4BX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.475 2.170 1.645 ;
        RECT  1.915 0.475 2.030 0.645 ;
        RECT  1.795 1.525 2.030 1.645 ;
        RECT  1.625 1.525 1.795 1.955 ;
        RECT  1.075 1.525 1.625 1.645 ;
        RECT  0.905 1.525 1.075 1.955 ;
        END
        AntennaDiffArea 0.643 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.770 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.010 1.200 1.270 ;
        RECT  0.910 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.410 1.005 1.610 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.235 1.375 ;
        END
        AntennaGateArea 0.0654 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.725 -0.210 2.240 0.210 ;
        RECT  0.555 -0.210 0.725 0.505 ;
        RECT  0.000 -0.210 0.555 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.155 2.310 2.240 2.730 ;
        RECT  1.985 1.845 2.155 2.730 ;
        RECT  1.435 2.310 1.985 2.730 ;
        RECT  1.265 1.845 1.435 2.730 ;
        RECT  0.715 2.310 1.265 2.730 ;
        RECT  0.545 1.845 0.715 2.730 ;
        RECT  0.000 2.310 0.545 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.790 0.765 1.910 1.270 ;
        RECT  1.720 0.765 1.790 0.885 ;
        RECT  1.600 0.625 1.720 0.885 ;
        RECT  0.510 0.625 1.600 0.745 ;
        RECT  0.390 0.625 0.510 1.625 ;
        RECT  0.335 0.625 0.390 0.745 ;
        RECT  0.335 1.505 0.390 1.625 ;
        RECT  0.165 0.565 0.335 0.745 ;
        RECT  0.165 1.505 0.335 1.675 ;
    END
END NAND4BX2AD
MACRO NAND4BX4AD
    CLASS CORE ;
    FOREIGN NAND4BX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.710 0.725 3.850 1.540 ;
        RECT  2.140 0.725 3.710 0.855 ;
        RECT  3.420 1.410 3.710 1.540 ;
        RECT  3.290 1.410 3.420 2.135 ;
        RECT  0.770 2.005 3.290 2.135 ;
        RECT  1.970 0.340 2.140 0.855 ;
        END
        AntennaDiffArea 1.206 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.210 1.020 3.330 1.280 ;
        RECT  3.170 1.160 3.210 1.280 ;
        RECT  3.050 1.160 3.170 1.885 ;
        RECT  0.910 1.765 3.050 1.885 ;
        RECT  0.790 1.685 0.910 1.885 ;
        RECT  0.770 1.685 0.790 1.805 ;
        RECT  0.630 1.040 0.770 1.805 ;
        END
        AntennaGateArea 0.3209 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.810 1.020 2.930 1.645 ;
        RECT  1.170 1.525 2.810 1.645 ;
        RECT  1.030 1.040 1.170 1.645 ;
        RECT  0.910 1.145 1.030 1.375 ;
        END
        AntennaGateArea 0.3226 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 1.000 2.570 1.405 ;
        RECT  1.610 1.285 2.450 1.405 ;
        RECT  1.390 1.040 1.610 1.405 ;
        END
        AntennaGateArea 0.3226 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.235 1.300 ;
        END
        AntennaGateArea 0.1295 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.545 -0.210 3.920 0.210 ;
        RECT  3.375 -0.210 3.545 0.550 ;
        RECT  0.690 -0.210 3.375 0.210 ;
        RECT  0.430 -0.210 0.690 0.505 ;
        RECT  0.000 -0.210 0.430 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.660 2.310 3.920 2.730 ;
        RECT  3.540 1.780 3.660 2.730 ;
        RECT  2.930 2.310 3.540 2.730 ;
        RECT  2.670 2.255 2.930 2.730 ;
        RECT  2.170 2.310 2.670 2.730 ;
        RECT  1.910 2.255 2.170 2.730 ;
        RECT  1.410 2.310 1.910 2.730 ;
        RECT  1.150 2.255 1.410 2.730 ;
        RECT  0.625 2.310 1.150 2.730 ;
        RECT  0.455 1.925 0.625 2.730 ;
        RECT  0.000 2.310 0.455 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  1.850 1.040 2.250 1.160 ;
        RECT  1.730 0.800 1.850 1.160 ;
        RECT  0.510 0.800 1.730 0.920 ;
        RECT  0.390 0.625 0.510 1.540 ;
        RECT  0.265 0.625 0.390 0.745 ;
        RECT  0.265 1.420 0.390 1.540 ;
        RECT  0.095 0.530 0.265 0.745 ;
        RECT  0.095 1.420 0.265 1.895 ;
    END
END NAND4BX4AD
MACRO NAND4BXLAD
    CLASS CORE ;
    FOREIGN NAND4BXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.565 2.170 1.615 ;
        RECT  1.915 0.565 2.030 0.735 ;
        RECT  1.735 1.495 2.030 1.615 ;
        RECT  1.565 1.495 1.735 1.680 ;
        RECT  1.015 1.495 1.565 1.615 ;
        RECT  0.845 1.495 1.015 1.680 ;
        END
        AntennaDiffArea 0.26 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 0.770 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.995 1.200 1.255 ;
        RECT  0.910 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 1.095 1.610 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.235 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.725 -0.210 2.240 0.210 ;
        RECT  0.555 -0.210 0.725 0.505 ;
        RECT  0.000 -0.210 0.555 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 2.310 2.240 2.730 ;
        RECT  1.880 1.735 2.140 2.730 ;
        RECT  1.420 2.310 1.880 2.730 ;
        RECT  1.160 1.735 1.420 2.730 ;
        RECT  0.700 2.310 1.160 2.730 ;
        RECT  0.440 1.735 0.700 2.730 ;
        RECT  0.000 2.310 0.440 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.760 0.855 1.880 1.130 ;
        RECT  1.720 0.855 1.760 0.975 ;
        RECT  1.600 0.625 1.720 0.975 ;
        RECT  0.510 0.625 1.600 0.745 ;
        RECT  0.390 0.625 0.510 1.615 ;
        RECT  0.335 0.625 0.390 0.745 ;
        RECT  0.275 1.495 0.390 1.615 ;
        RECT  0.165 0.565 0.335 0.745 ;
        RECT  0.105 1.495 0.275 1.680 ;
    END
END NAND4BXLAD
MACRO NAND4X1AD
    CLASS CORE ;
    FOREIGN NAND4X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.490 0.525 1.610 1.620 ;
        RECT  1.450 0.525 1.490 0.815 ;
        RECT  1.275 1.500 1.490 1.620 ;
        RECT  1.105 1.500 1.275 2.005 ;
        RECT  0.575 1.500 1.105 1.620 ;
        RECT  0.405 1.500 0.575 2.005 ;
        END
        AntennaDiffArea 0.383 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.230 1.375 ;
        END
        AntennaGateArea 0.0904 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.010 0.700 1.270 ;
        RECT  0.350 0.865 0.490 1.375 ;
        END
        AntennaGateArea 0.0904 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.865 1.070 1.375 ;
        END
        AntennaGateArea 0.0904 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 0.980 1.370 1.240 ;
        RECT  1.190 0.865 1.330 1.375 ;
        END
        AntennaGateArea 0.0904 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.255 -0.210 1.680 0.210 ;
        RECT  0.085 -0.210 0.255 0.725 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.565 2.310 1.680 2.730 ;
        RECT  1.395 2.265 1.565 2.730 ;
        RECT  0.925 2.310 1.395 2.730 ;
        RECT  0.755 2.265 0.925 2.730 ;
        RECT  0.285 2.310 0.755 2.730 ;
        RECT  0.115 2.265 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
	 END
END NAND4X1AD
MACRO NAND4X2AD
    CLASS CORE ;
    FOREIGN NAND4X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.585 1.890 1.620 ;
        RECT  1.750 0.365 1.760 1.620 ;
        RECT  1.500 0.365 1.750 0.745 ;
        RECT  1.415 1.500 1.750 1.620 ;
        RECT  1.245 1.500 1.415 2.005 ;
        RECT  0.695 1.500 1.245 1.620 ;
        RECT  0.525 1.500 0.695 2.005 ;
        END
        AntennaDiffArea 0.671 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.310 0.845 0.490 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 0.865 0.790 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.080 1.020 1.180 1.280 ;
        RECT  0.910 0.865 1.080 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.865 1.610 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.365 -0.210 1.960 0.210 ;
        RECT  0.195 -0.210 0.365 0.675 ;
        RECT  0.000 -0.210 0.195 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.775 2.310 1.960 2.730 ;
        RECT  1.605 1.740 1.775 2.730 ;
        RECT  1.055 2.310 1.605 2.730 ;
        RECT  0.885 1.740 1.055 2.730 ;
        RECT  0.305 2.310 0.885 2.730 ;
        RECT  0.135 1.585 0.305 2.730 ;
        RECT  0.000 2.310 0.135 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
	 END
END NAND4X2AD
MACRO NAND4X4AD
    CLASS CORE ;
    FOREIGN NAND4X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.145 0.770 3.290 2.010 ;
        RECT  2.765 0.770 3.145 0.900 ;
        RECT  0.400 1.880 3.145 2.010 ;
        RECT  2.635 0.380 2.765 0.900 ;
        RECT  1.435 0.380 2.635 0.500 ;
        END
        AntennaDiffArea 1.21 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.020 2.840 1.760 ;
        RECT  0.510 1.640 2.720 1.760 ;
        RECT  0.390 1.500 0.510 1.760 ;
        RECT  0.235 1.500 0.390 1.655 ;
        RECT  0.070 1.020 0.235 1.655 ;
        END
        AntennaGateArea 0.324 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.370 1.020 2.495 1.520 ;
        RECT  0.770 1.400 2.370 1.520 ;
        RECT  0.630 0.865 0.770 1.520 ;
        RECT  0.560 1.020 0.630 1.280 ;
        END
        AntennaGateArea 0.324 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.060 0.620 2.180 1.260 ;
        RECT  1.050 0.620 2.060 0.740 ;
        RECT  0.910 0.585 1.050 1.260 ;
        END
        AntennaGateArea 0.324 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.040 1.790 1.160 ;
        RECT  1.190 0.865 1.330 1.160 ;
        END
        AntennaGateArea 0.324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.200 -0.210 3.360 0.210 ;
        RECT  2.940 -0.210 3.200 0.650 ;
        RECT  0.255 -0.210 2.940 0.210 ;
        RECT  0.085 -0.210 0.255 0.785 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.180 2.310 3.360 2.730 ;
        RECT  2.920 2.130 3.180 2.730 ;
        RECT  2.460 2.310 2.920 2.730 ;
        RECT  2.200 2.130 2.460 2.730 ;
        RECT  1.740 2.310 2.200 2.730 ;
        RECT  1.480 2.130 1.740 2.730 ;
        RECT  1.020 2.310 1.480 2.730 ;
        RECT  0.760 2.130 1.020 2.730 ;
        RECT  0.255 2.310 0.760 2.730 ;
        RECT  0.085 1.845 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
	 END
END NAND4X4AD
MACRO NAND4X6AD
    CLASS CORE ;
    FOREIGN NAND4X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.800 0.685 4.970 1.665 ;
        RECT  4.730 0.685 4.800 0.855 ;
        RECT  4.465 1.485 4.800 1.665 ;
        RECT  4.560 0.380 4.730 0.855 ;
        RECT  4.295 1.485 4.465 1.940 ;
        RECT  3.705 1.485 4.295 1.665 ;
        RECT  3.535 1.485 3.705 1.935 ;
        RECT  3.210 1.485 3.535 1.665 ;
        RECT  3.045 1.485 3.210 2.100 ;
        RECT  3.040 1.485 3.045 2.140 ;
        RECT  0.230 1.980 3.040 2.140 ;
        RECT  1.560 0.360 1.730 0.790 ;
        RECT  0.230 0.535 1.560 0.705 ;
        RECT  0.070 0.535 0.230 2.140 ;
        END
        AntennaDiffArea 1.826 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.920 1.140 3.390 1.260 ;
        RECT  2.800 1.140 2.920 1.860 ;
        RECT  0.490 1.740 2.800 1.860 ;
        RECT  0.350 1.020 0.490 1.860 ;
        END
        AntennaGateArea 0.4812 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.710 0.895 3.830 1.280 ;
        RECT  2.620 0.895 3.710 1.020 ;
        RECT  2.500 0.895 2.620 1.620 ;
        RECT  0.770 1.500 2.500 1.620 ;
        RECT  0.630 0.865 0.770 1.620 ;
        END
        AntennaGateArea 0.4808 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.080 0.655 4.200 1.280 ;
        RECT  2.290 0.655 4.080 0.775 ;
        RECT  2.170 0.655 2.290 1.380 ;
        RECT  1.190 1.260 2.170 1.380 ;
        RECT  1.050 1.120 1.190 1.380 ;
        RECT  0.910 0.865 1.050 1.380 ;
        END
        AntennaGateArea 0.4808 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.440 1.020 4.530 1.280 ;
        RECT  4.320 0.415 4.440 1.280 ;
        RECT  2.020 0.415 4.320 0.535 ;
        RECT  1.900 0.415 2.020 1.140 ;
        RECT  1.705 0.910 1.900 1.140 ;
        RECT  1.425 1.020 1.705 1.140 ;
        END
        AntennaGateArea 0.4808 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.310 -0.210 5.040 0.210 ;
        RECT  3.050 -0.210 3.310 0.290 ;
        RECT  0.255 -0.210 3.050 0.210 ;
        RECT  0.085 -0.210 0.255 0.415 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.825 2.310 5.040 2.730 ;
        RECT  4.655 1.825 4.825 2.730 ;
        RECT  4.085 2.310 4.655 2.730 ;
        RECT  3.915 1.825 4.085 2.730 ;
        RECT  3.370 2.310 3.915 2.730 ;
        RECT  3.110 2.280 3.370 2.730 ;
        RECT  2.610 2.310 3.110 2.730 ;
        RECT  2.350 2.280 2.610 2.730 ;
        RECT  1.850 2.310 2.350 2.730 ;
        RECT  1.590 2.280 1.850 2.730 ;
        RECT  1.090 2.310 1.590 2.730 ;
        RECT  0.830 2.280 1.090 2.730 ;
        RECT  0.330 2.310 0.830 2.730 ;
        RECT  0.070 2.280 0.330 2.730 ;
        RECT  0.000 2.310 0.070 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.040 2.520 ;
	 END
END NAND4X6AD
MACRO NAND4X8AD
    CLASS CORE ;
    FOREIGN NAND4X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.220 0.600 6.470 2.140 ;
        RECT  5.715 0.600 6.220 0.850 ;
        RECT  0.230 1.980 6.220 2.140 ;
        RECT  5.205 0.490 5.715 0.910 ;
        RECT  4.850 0.600 5.205 0.850 ;
        RECT  4.610 0.360 4.850 0.850 ;
        RECT  1.560 0.360 1.730 0.790 ;
        RECT  0.230 0.535 1.560 0.745 ;
        RECT  0.070 0.535 0.230 2.140 ;
        END
        AntennaDiffArea 2.412 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.930 1.020 6.050 1.860 ;
        RECT  3.480 1.740 5.930 1.860 ;
        RECT  3.360 1.140 3.480 1.860 ;
        RECT  2.920 1.140 3.360 1.260 ;
        RECT  2.800 1.140 2.920 1.860 ;
        RECT  0.490 1.740 2.800 1.860 ;
        RECT  0.350 1.020 0.490 1.860 ;
        END
        AntennaGateArea 0.6416 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.660 1.090 5.800 1.210 ;
        RECT  5.540 1.090 5.660 1.620 ;
        RECT  3.830 1.500 5.540 1.620 ;
        RECT  3.710 0.895 3.830 1.620 ;
        RECT  2.620 0.895 3.710 1.020 ;
        RECT  2.500 0.895 2.620 1.620 ;
        RECT  0.770 1.500 2.500 1.620 ;
        RECT  0.630 0.865 0.770 1.620 ;
        END
        AntennaGateArea 0.6416 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.300 1.090 5.420 1.210 ;
        RECT  5.160 1.090 5.300 1.380 ;
        RECT  4.200 1.260 5.160 1.380 ;
        RECT  4.080 0.655 4.200 1.380 ;
        RECT  2.290 0.655 4.080 0.775 ;
        RECT  2.170 0.655 2.290 1.380 ;
        RECT  1.190 1.260 2.170 1.380 ;
        RECT  1.050 1.120 1.190 1.380 ;
        RECT  0.910 0.865 1.050 1.380 ;
        END
        AntennaGateArea 0.6416 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.440 1.020 4.890 1.140 ;
        RECT  4.320 0.415 4.440 1.140 ;
        RECT  2.020 0.415 4.320 0.535 ;
        RECT  1.900 0.415 2.020 1.140 ;
        RECT  1.705 0.910 1.900 1.140 ;
        RECT  1.425 1.020 1.705 1.140 ;
        END
        AntennaGateArea 0.6416 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.225 -0.210 6.720 0.210 ;
        RECT  6.055 -0.210 6.225 0.415 ;
        RECT  3.310 -0.210 6.055 0.210 ;
        RECT  3.050 -0.210 3.310 0.290 ;
        RECT  0.255 -0.210 3.050 0.210 ;
        RECT  0.085 -0.210 0.255 0.415 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.410 2.310 6.720 2.730 ;
        RECT  6.150 2.280 6.410 2.730 ;
        RECT  5.650 2.310 6.150 2.730 ;
        RECT  5.390 2.280 5.650 2.730 ;
        RECT  4.890 2.310 5.390 2.730 ;
        RECT  4.630 2.280 4.890 2.730 ;
        RECT  4.130 2.310 4.630 2.730 ;
        RECT  3.870 2.280 4.130 2.730 ;
        RECT  3.370 2.310 3.870 2.730 ;
        RECT  3.110 2.280 3.370 2.730 ;
        RECT  2.610 2.310 3.110 2.730 ;
        RECT  2.350 2.280 2.610 2.730 ;
        RECT  1.850 2.310 2.350 2.730 ;
        RECT  1.590 2.280 1.850 2.730 ;
        RECT  1.090 2.310 1.590 2.730 ;
        RECT  0.830 2.280 1.090 2.730 ;
        RECT  0.330 2.310 0.830 2.730 ;
        RECT  0.070 2.280 0.330 2.730 ;
        RECT  0.000 2.310 0.070 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.720 2.520 ;
	 END
END NAND4X8AD
MACRO NAND4XLAD
    CLASS CORE ;
    FOREIGN NAND4XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.490 0.510 1.610 1.620 ;
        RECT  1.450 0.510 1.490 0.815 ;
        RECT  1.275 1.500 1.490 1.620 ;
        RECT  1.105 1.500 1.275 1.670 ;
        RECT  0.575 1.500 1.105 1.620 ;
        RECT  0.405 1.500 0.575 1.670 ;
        END
        AntennaDiffArea 0.254 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.230 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.010 0.700 1.270 ;
        RECT  0.350 0.865 0.490 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.865 1.070 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 0.980 1.370 1.240 ;
        RECT  1.190 0.865 1.330 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.255 -0.210 1.680 0.210 ;
        RECT  0.085 -0.210 0.255 0.725 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.565 2.310 1.680 2.730 ;
        RECT  1.395 2.055 1.565 2.730 ;
        RECT  0.925 2.310 1.395 2.730 ;
        RECT  0.755 2.055 0.925 2.730 ;
        RECT  0.285 2.310 0.755 2.730 ;
        RECT  0.115 2.055 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
	 END
END NAND4XLAD
MACRO NOR2BX1AD
    CLASS CORE ;
    FOREIGN NOR2BX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.185 0.670 1.330 1.860 ;
        RECT  0.755 0.670 1.185 0.820 ;
        RECT  1.160 1.340 1.185 1.860 ;
        END
        AntennaDiffArea 0.222 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.000 0.800 1.655 ;
        END
        AntennaGateArea 0.0904 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.010 0.490 1.655 ;
        END
        AntennaGateArea 0.0424 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.175 -0.210 1.400 0.210 ;
        RECT  0.485 -0.210 1.175 0.380 ;
        RECT  0.000 -0.210 0.485 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.710 2.310 1.400 2.730 ;
        RECT  0.450 2.015 0.710 2.730 ;
        RECT  0.000 2.310 0.450 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.990 2.070 1.230 2.190 ;
        RECT  0.870 1.775 0.990 2.190 ;
        RECT  0.230 1.775 0.870 1.895 ;
        RECT  0.190 0.730 0.265 0.900 ;
        RECT  0.190 1.340 0.230 1.895 ;
        RECT  0.070 0.730 0.190 1.895 ;
    END
END NOR2BX1AD
MACRO NOR2BX2AD
    CLASS CORE ;
    FOREIGN NOR2BX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.735 1.610 1.950 ;
        RECT  1.105 0.735 1.470 0.875 ;
        RECT  1.465 1.735 1.470 1.950 ;
        RECT  1.295 1.735 1.465 2.165 ;
        RECT  0.935 0.355 1.105 0.875 ;
        END
        AntennaDiffArea 0.394 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.010 1.050 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.015 0.595 1.375 ;
        END
        AntennaGateArea 0.0652 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.465 -0.210 1.680 0.210 ;
        RECT  1.295 -0.210 1.465 0.615 ;
        RECT  0.745 -0.210 1.295 0.210 ;
        RECT  0.575 -0.210 0.745 0.785 ;
        RECT  0.000 -0.210 0.575 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.835 2.310 1.680 2.730 ;
        RECT  0.665 1.735 0.835 2.730 ;
        RECT  0.000 2.310 0.665 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.290 1.055 1.345 1.225 ;
        RECT  1.170 1.055 1.290 1.615 ;
        RECT  0.230 1.495 1.170 1.615 ;
        RECT  0.230 0.695 0.365 0.865 ;
        RECT  0.110 0.695 0.230 1.615 ;
    END
END NOR2BX2AD
MACRO NOR2BX4AD
    CLASS CORE ;
    FOREIGN NOR2BX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.795 2.170 1.605 ;
        RECT  1.770 0.795 2.030 0.915 ;
        RECT  1.350 1.465 2.030 1.605 ;
        RECT  1.650 0.330 1.770 0.915 ;
        RECT  1.600 0.330 1.650 0.760 ;
        RECT  1.045 0.640 1.600 0.760 ;
        RECT  1.180 1.465 1.350 2.155 ;
        RECT  0.875 0.330 1.045 0.760 ;
        END
        AntennaDiffArea 0.71 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.655 1.065 1.895 1.235 ;
        RECT  1.515 1.065 1.655 1.330 ;
        RECT  1.395 0.880 1.515 1.330 ;
        RECT  0.800 0.880 1.395 1.000 ;
        RECT  0.680 0.880 0.800 1.270 ;
        END
        AntennaGateArea 0.324 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.510 1.285 ;
        RECT  0.325 1.010 0.350 1.285 ;
        END
        AntennaGateArea 0.129 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.135 -0.210 2.240 0.210 ;
        RECT  1.965 -0.210 2.135 0.675 ;
        RECT  1.405 -0.210 1.965 0.210 ;
        RECT  1.235 -0.210 1.405 0.520 ;
        RECT  0.685 -0.210 1.235 0.210 ;
        RECT  0.515 -0.210 0.685 0.715 ;
        RECT  0.000 -0.210 0.515 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.015 2.310 2.240 2.730 ;
        RECT  1.845 1.725 2.015 2.730 ;
        RECT  0.685 2.310 1.845 2.730 ;
        RECT  0.515 1.655 0.685 2.730 ;
        RECT  0.000 2.310 0.515 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.040 1.120 1.275 1.240 ;
        RECT  0.920 1.120 1.040 1.535 ;
        RECT  0.325 1.415 0.920 1.535 ;
        RECT  0.205 0.330 0.370 0.720 ;
        RECT  0.205 1.415 0.325 1.950 ;
        RECT  0.155 0.330 0.205 1.950 ;
        RECT  0.110 0.330 0.155 1.535 ;
        RECT  0.085 0.520 0.110 1.535 ;
    END
END NOR2BX4AD
MACRO NOR2BX8AD
    CLASS CORE ;
    FOREIGN NOR2BX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.860 0.540 4.100 1.820 ;
        RECT  3.705 0.540 3.860 0.710 ;
        RECT  3.475 1.580 3.860 1.820 ;
        RECT  3.445 0.330 3.705 0.710 ;
        RECT  2.965 1.580 3.475 2.030 ;
        RECT  2.945 0.540 3.445 0.710 ;
        RECT  1.760 1.580 2.965 1.820 ;
        RECT  2.685 0.330 2.945 0.710 ;
        RECT  2.185 0.540 2.685 0.710 ;
        RECT  1.925 0.330 2.185 0.710 ;
        RECT  1.425 0.540 1.925 0.710 ;
        RECT  1.590 1.465 1.760 2.155 ;
        RECT  1.165 0.330 1.425 0.710 ;
        END
        AntennaDiffArea 1.242 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.615 0.880 3.735 1.295 ;
        RECT  2.780 0.880 3.615 1.000 ;
        RECT  2.260 0.880 2.780 1.170 ;
        RECT  1.205 0.880 2.260 1.000 ;
        RECT  1.085 0.880 1.205 1.280 ;
        END
        AntennaGateArea 0.648 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.205 1.085 0.725 1.330 ;
        END
        AntennaGateArea 0.2619 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.045 -0.210 4.200 0.210 ;
        RECT  3.875 -0.210 4.045 0.420 ;
        RECT  3.280 -0.210 3.875 0.210 ;
        RECT  3.110 -0.210 3.280 0.420 ;
        RECT  2.520 -0.210 3.110 0.210 ;
        RECT  2.350 -0.210 2.520 0.420 ;
        RECT  1.760 -0.210 2.350 0.210 ;
        RECT  1.590 -0.210 1.760 0.420 ;
        RECT  1.000 -0.210 1.590 0.210 ;
        RECT  0.830 -0.210 1.000 0.725 ;
        RECT  0.265 -0.210 0.830 0.210 ;
        RECT  0.095 -0.210 0.265 0.860 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.910 2.310 4.200 2.730 ;
        RECT  3.740 1.940 3.910 2.730 ;
        RECT  2.555 2.310 3.740 2.730 ;
        RECT  2.385 1.940 2.555 2.730 ;
        RECT  1.020 2.310 2.385 2.730 ;
        RECT  0.850 1.735 1.020 2.730 ;
        RECT  0.265 2.310 0.850 2.730 ;
        RECT  0.095 1.525 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  3.065 1.125 3.465 1.245 ;
        RECT  2.945 1.125 3.065 1.410 ;
        RECT  2.105 1.290 2.945 1.410 ;
        RECT  1.985 1.120 2.105 1.410 ;
        RECT  1.445 1.120 1.985 1.240 ;
        RECT  1.325 1.120 1.445 1.600 ;
        RECT  0.965 1.480 1.325 1.600 ;
        RECT  0.845 0.845 0.965 1.600 ;
        RECT  0.625 0.845 0.845 0.965 ;
        RECT  0.625 1.480 0.845 1.600 ;
        RECT  0.455 0.430 0.625 0.965 ;
        RECT  0.455 1.480 0.625 1.955 ;
    END
END NOR2BX8AD
MACRO NOR2BXLAD
    CLASS CORE ;
    FOREIGN NOR2BXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.210 0.755 1.330 1.675 ;
        RECT  0.760 0.755 1.210 0.875 ;
        RECT  1.160 1.415 1.210 1.675 ;
        END
        AntennaDiffArea 0.144 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.000 0.800 1.655 ;
        END
        AntennaGateArea 0.0604 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.010 0.490 1.655 ;
        END
        AntennaGateArea 0.0404 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.175 -0.210 1.400 0.210 ;
        RECT  0.485 -0.210 1.175 0.380 ;
        RECT  0.000 -0.210 0.485 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.710 2.310 1.400 2.730 ;
        RECT  0.450 2.015 0.710 2.730 ;
        RECT  0.000 2.310 0.450 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.990 1.880 1.230 2.000 ;
        RECT  0.870 1.775 0.990 2.000 ;
        RECT  0.230 1.775 0.870 1.895 ;
        RECT  0.190 0.730 0.265 0.900 ;
        RECT  0.190 1.330 0.230 1.895 ;
        RECT  0.070 0.730 0.190 1.895 ;
    END
END NOR2BXLAD
MACRO NOR2X1AD
    CLASS CORE ;
    FOREIGN NOR2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.700 1.050 1.655 ;
        RECT  0.440 0.700 0.910 0.840 ;
        RECT  0.905 1.495 0.910 1.655 ;
        RECT  0.735 1.495 0.905 1.925 ;
        END
        AntennaDiffArea 0.216 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.000 0.490 1.655 ;
        RECT  0.260 1.000 0.350 1.265 ;
        END
        AntennaGateArea 0.09 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 0.990 0.780 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.035 -0.210 1.120 0.210 ;
        RECT  0.865 -0.210 1.035 0.580 ;
        RECT  0.290 -0.210 0.865 0.210 ;
        RECT  0.130 -0.210 0.290 0.880 ;
        RECT  0.000 -0.210 0.130 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.230 2.310 1.120 2.730 ;
        RECT  0.090 1.410 0.230 2.730 ;
        RECT  0.000 2.310 0.090 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
	 END
END NOR2X1AD
MACRO NOR2X2AD
    CLASS CORE ;
    FOREIGN NOR2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.000 0.730 1.050 1.935 ;
        RECT  0.910 0.730 1.000 2.175 ;
        RECT  0.625 0.730 0.910 0.875 ;
        RECT  0.740 1.795 0.910 2.175 ;
        RECT  0.455 0.360 0.625 0.875 ;
        END
        AntennaDiffArea 0.394 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.010 0.490 1.375 ;
        RECT  0.070 1.140 0.330 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.010 0.780 1.655 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.985 -0.210 1.120 0.210 ;
        RECT  0.815 -0.210 0.985 0.610 ;
        RECT  0.265 -0.210 0.815 0.210 ;
        RECT  0.095 -0.210 0.265 0.790 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.345 2.310 1.120 2.730 ;
        RECT  0.175 1.605 0.345 2.730 ;
        RECT  0.000 2.310 0.175 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
	 END
END NOR2X2AD
MACRO NOR2X3AD
    CLASS CORE ;
    FOREIGN NOR2X3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.625 1.810 1.610 ;
        RECT  0.450 0.625 1.670 0.765 ;
        RECT  1.055 1.470 1.670 1.610 ;
        RECT  0.885 1.470 1.055 1.900 ;
        END
        AntennaDiffArea 0.494 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.355 0.890 1.550 1.315 ;
        RECT  0.535 0.890 1.355 1.010 ;
        RECT  0.305 0.890 0.535 1.285 ;
        END
        AntennaGateArea 0.2445 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.130 1.230 1.330 ;
        END
        AntennaGateArea 0.245 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.825 -0.210 1.960 0.210 ;
        RECT  1.655 -0.210 1.825 0.505 ;
        RECT  1.055 -0.210 1.655 0.210 ;
        RECT  0.885 -0.210 1.055 0.505 ;
        RECT  0.300 -0.210 0.885 0.210 ;
        RECT  0.130 -0.210 0.300 0.735 ;
        RECT  0.000 -0.210 0.130 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.685 2.310 1.960 2.730 ;
        RECT  1.515 1.730 1.685 2.730 ;
        RECT  0.415 2.310 1.515 2.730 ;
        RECT  0.245 1.470 0.415 2.730 ;
        RECT  0.000 2.310 0.245 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
	 END
END NOR2X3AD
MACRO NOR2X4AD
    CLASS CORE ;
    FOREIGN NOR2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.780 1.890 1.760 ;
        RECT  1.400 0.780 1.750 0.920 ;
        RECT  1.040 1.620 1.750 1.760 ;
        RECT  1.230 0.340 1.400 0.920 ;
        RECT  0.725 0.605 1.230 0.745 ;
        RECT  0.870 1.620 1.040 2.050 ;
        RECT  0.465 0.365 0.725 0.745 ;
        END
        AntennaDiffArea 0.602 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.395 1.040 1.515 1.500 ;
        RECT  0.510 1.380 1.395 1.500 ;
        RECT  0.350 1.000 0.510 1.500 ;
        END
        AntennaGateArea 0.3249 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.000 1.130 1.260 ;
        RECT  0.630 0.865 1.050 1.260 ;
        END
        AntennaGateArea 0.324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.805 -0.210 1.960 0.210 ;
        RECT  1.545 -0.210 1.805 0.660 ;
        RECT  1.040 -0.210 1.545 0.210 ;
        RECT  0.870 -0.210 1.040 0.485 ;
        RECT  0.320 -0.210 0.870 0.210 ;
        RECT  0.150 -0.210 0.320 0.795 ;
        RECT  0.000 -0.210 0.150 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.650 2.310 1.960 2.730 ;
        RECT  1.480 1.880 1.650 2.730 ;
        RECT  0.430 2.310 1.480 2.730 ;
        RECT  0.260 1.620 0.430 2.730 ;
        RECT  0.000 2.310 0.260 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
	 END
END NOR2X4AD
MACRO NOR2X5AD
    CLASS CORE ;
    FOREIGN NOR2X5AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.340 0.730 2.450 1.795 ;
        RECT  2.310 0.730 2.340 2.105 ;
        RECT  2.070 0.730 2.310 0.870 ;
        RECT  2.170 1.570 2.310 2.105 ;
        RECT  1.015 1.570 2.170 1.710 ;
        RECT  1.900 0.420 2.070 0.870 ;
        RECT  1.350 0.730 1.900 0.870 ;
        RECT  1.180 0.425 1.350 0.870 ;
        RECT  0.630 0.730 1.180 0.870 ;
        RECT  0.845 1.570 1.015 2.105 ;
        RECT  0.460 0.420 0.630 0.870 ;
        END
        AntennaDiffArea 0.855 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.495 1.010 1.845 1.150 ;
        RECT  0.490 1.010 0.495 1.270 ;
        RECT  0.255 1.010 0.490 1.375 ;
        END
        AntennaGateArea 0.402 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.115 2.170 1.430 ;
        RECT  0.680 1.290 2.030 1.430 ;
        END
        AntennaGateArea 0.402 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 -0.210 2.520 0.210 ;
        RECT  2.260 -0.210 2.430 0.605 ;
        RECT  1.710 -0.210 2.260 0.210 ;
        RECT  1.540 -0.210 1.710 0.605 ;
        RECT  0.990 -0.210 1.540 0.210 ;
        RECT  0.820 -0.210 0.990 0.605 ;
        RECT  0.270 -0.210 0.820 0.210 ;
        RECT  0.100 -0.210 0.270 0.850 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.685 2.310 2.520 2.730 ;
        RECT  1.515 1.845 1.685 2.730 ;
        RECT  0.370 2.310 1.515 2.730 ;
        RECT  0.200 1.585 0.370 2.730 ;
        RECT  0.000 2.310 0.200 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
	 END
END NOR2X5AD
MACRO NOR2X6AD
    CLASS CORE ;
    FOREIGN NOR2X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.305 0.605 2.450 1.730 ;
        RECT  2.280 0.605 2.305 2.040 ;
        RECT  2.055 0.605 2.280 0.775 ;
        RECT  2.135 1.560 2.280 2.040 ;
        RECT  0.990 1.560 2.135 1.730 ;
        RECT  1.885 0.345 2.055 0.775 ;
        RECT  1.335 0.605 1.885 0.775 ;
        RECT  1.165 0.345 1.335 0.775 ;
        RECT  0.615 0.605 1.165 0.775 ;
        RECT  0.820 1.560 0.990 2.040 ;
        RECT  0.445 0.345 0.615 0.775 ;
        END
        AntennaDiffArea 1.024 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.135 1.610 1.440 ;
        RECT  0.460 1.315 1.350 1.440 ;
        RECT  0.340 1.020 0.460 1.440 ;
        END
        AntennaGateArea 0.486 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.895 2.130 1.275 ;
        RECT  1.160 0.895 2.010 1.015 ;
        RECT  0.690 0.895 1.160 1.195 ;
        END
        AntennaGateArea 0.486 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.415 -0.210 2.520 0.210 ;
        RECT  2.245 -0.210 2.415 0.485 ;
        RECT  1.695 -0.210 2.245 0.210 ;
        RECT  1.525 -0.210 1.695 0.485 ;
        RECT  0.975 -0.210 1.525 0.210 ;
        RECT  0.805 -0.210 0.975 0.485 ;
        RECT  0.255 -0.210 0.805 0.210 ;
        RECT  0.085 -0.210 0.255 0.775 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.655 2.310 2.520 2.730 ;
        RECT  1.485 1.850 1.655 2.730 ;
        RECT  0.365 2.310 1.485 2.730 ;
        RECT  0.195 1.610 0.365 2.730 ;
        RECT  0.000 2.310 0.195 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
	 END
END NOR2X6AD
MACRO NOR2X8AD
    CLASS CORE ;
    FOREIGN NOR2X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.615 0.335 2.785 0.765 ;
        RECT  2.125 1.585 2.635 2.030 ;
        RECT  2.065 0.595 2.615 0.765 ;
        RECT  0.995 1.585 2.125 1.835 ;
        RECT  1.895 0.335 2.065 0.765 ;
        RECT  1.345 0.595 1.895 0.765 ;
        RECT  1.175 0.335 1.345 0.765 ;
        RECT  0.625 0.595 1.175 0.765 ;
        RECT  0.825 1.585 0.995 2.015 ;
        RECT  0.260 1.585 0.825 1.835 ;
        RECT  0.455 0.335 0.625 0.765 ;
        RECT  0.260 0.595 0.455 0.765 ;
        RECT  0.090 0.595 0.260 1.835 ;
        END
        AntennaDiffArea 1.334 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.770 0.885 2.890 1.270 ;
        RECT  1.845 0.885 2.770 1.005 ;
        RECT  1.325 0.885 1.845 1.175 ;
        RECT  0.500 0.885 1.325 1.005 ;
        RECT  0.380 0.885 0.500 1.280 ;
        END
        AntennaGateArea 0.648 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.125 2.500 1.245 ;
        RECT  1.980 1.125 2.170 1.415 ;
        RECT  1.170 1.295 1.980 1.415 ;
        RECT  1.030 1.125 1.170 1.415 ;
        RECT  0.650 1.125 1.030 1.245 ;
        END
        AntennaGateArea 0.648 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.145 -0.210 3.360 0.210 ;
        RECT  2.975 -0.210 3.145 0.765 ;
        RECT  2.425 -0.210 2.975 0.210 ;
        RECT  2.255 -0.210 2.425 0.475 ;
        RECT  1.705 -0.210 2.255 0.210 ;
        RECT  1.535 -0.210 1.705 0.475 ;
        RECT  0.985 -0.210 1.535 0.210 ;
        RECT  0.815 -0.210 0.985 0.475 ;
        RECT  0.265 -0.210 0.815 0.210 ;
        RECT  0.095 -0.210 0.265 0.475 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.040 2.310 3.360 2.730 ;
        RECT  2.870 1.485 3.040 2.730 ;
        RECT  1.665 2.310 2.870 2.730 ;
        RECT  1.495 1.955 1.665 2.730 ;
        RECT  0.375 2.310 1.495 2.730 ;
        RECT  0.205 1.955 0.375 2.730 ;
        RECT  0.000 2.310 0.205 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
	 END
END NOR2X8AD
MACRO NOR2XLAD
    CLASS CORE ;
    FOREIGN NOR2XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.750 1.050 1.670 ;
        RECT  0.410 0.750 0.910 0.890 ;
        RECT  0.705 1.500 0.910 1.670 ;
        END
        AntennaDiffArea 0.144 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.025 0.490 1.655 ;
        RECT  0.270 1.025 0.350 1.285 ;
        END
        AntennaGateArea 0.06 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.010 0.790 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.005 -0.210 1.120 0.210 ;
        RECT  0.835 -0.210 1.005 0.630 ;
        RECT  0.265 -0.210 0.835 0.210 ;
        RECT  0.095 -0.210 0.265 0.905 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.230 2.310 1.120 2.730 ;
        RECT  0.110 1.455 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.120 2.520 ;
	 END
END NOR2XLAD
MACRO NOR3BX1AD
    CLASS CORE ;
    FOREIGN NOR3BX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.690 1.610 1.925 ;
        RECT  1.425 0.690 1.470 0.860 ;
        RECT  1.445 1.405 1.470 1.925 ;
        RECT  0.925 0.740 1.425 0.860 ;
        RECT  0.755 0.690 0.925 0.860 ;
        END
        AntennaDiffArea 0.283 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.000 0.770 1.420 ;
        END
        AntennaGateArea 0.0904 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.015 1.065 1.415 ;
        END
        AntennaGateArea 0.09 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.010 0.270 1.270 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.0424 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.185 -0.210 1.680 0.210 ;
        RECT  0.495 -0.210 1.185 0.325 ;
        RECT  0.000 -0.210 0.495 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.605 2.310 1.680 2.730 ;
        RECT  0.435 1.935 0.605 2.730 ;
        RECT  0.000 2.310 0.435 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.305 1.020 1.350 1.280 ;
        RECT  1.185 1.020 1.305 1.665 ;
        RECT  0.510 1.545 1.185 1.665 ;
        RECT  0.390 0.625 0.510 1.665 ;
        RECT  0.330 0.625 0.390 0.745 ;
        RECT  0.085 1.495 0.390 1.665 ;
        RECT  0.210 0.330 0.330 0.745 ;
        RECT  0.070 0.330 0.210 0.450 ;
    END
END NOR3BX1AD
MACRO NOR3BX2AD
    CLASS CORE ;
    FOREIGN NOR3BX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 0.605 1.890 1.960 ;
        RECT  1.755 0.330 1.800 1.960 ;
        RECT  1.750 0.330 1.755 2.170 ;
        RECT  1.540 0.330 1.750 0.745 ;
        RECT  1.585 1.740 1.750 2.170 ;
        RECT  1.080 0.605 1.540 0.745 ;
        RECT  0.820 0.330 1.080 0.745 ;
        END
        AntennaDiffArea 0.553 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.010 0.860 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.865 1.330 1.280 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.990 0.510 1.375 ;
        END
        AntennaGateArea 0.0651 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.395 -0.210 1.960 0.210 ;
        RECT  1.225 -0.210 1.395 0.485 ;
        RECT  0.675 -0.210 1.225 0.210 ;
        RECT  0.505 -0.210 0.675 0.745 ;
        RECT  0.000 -0.210 0.505 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.795 2.310 1.960 2.730 ;
        RECT  0.625 1.740 0.795 2.730 ;
        RECT  0.000 2.310 0.625 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.460 1.010 1.580 1.620 ;
        RECT  0.230 1.500 1.460 1.620 ;
        RECT  0.230 0.700 0.295 0.870 ;
        RECT  0.110 0.700 0.230 1.620 ;
    END
END NOR3BX2AD
MACRO NOR3BX4AD
    CLASS CORE ;
    FOREIGN NOR3BX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 0.825 3.010 1.940 ;
        RECT  2.560 0.825 2.870 0.965 ;
        RECT  1.870 1.800 2.870 1.940 ;
        RECT  2.320 0.370 2.560 0.965 ;
        RECT  2.300 0.370 2.320 0.780 ;
        RECT  1.840 0.640 2.300 0.780 ;
        RECT  1.610 1.800 1.870 2.190 ;
        RECT  1.580 0.370 1.840 0.780 ;
        RECT  1.120 0.640 1.580 0.780 ;
        RECT  0.860 0.370 1.120 0.780 ;
        END
        AntennaDiffArea 0.838 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.085 2.695 1.255 ;
        RECT  2.470 1.085 2.590 1.680 ;
        RECT  1.095 1.560 2.470 1.680 ;
        RECT  0.980 1.470 1.095 1.680 ;
        RECT  0.860 1.140 0.980 1.680 ;
        RECT  0.720 1.140 0.860 1.260 ;
        END
        AntennaGateArea 0.3249 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.085 2.335 1.255 ;
        RECT  2.030 1.085 2.170 1.440 ;
        RECT  1.395 1.320 2.030 1.440 ;
        RECT  1.275 1.140 1.395 1.440 ;
        RECT  1.100 1.140 1.275 1.260 ;
        END
        AntennaGateArea 0.3259 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.100 1.025 0.360 1.375 ;
        RECT  0.070 1.140 0.100 1.375 ;
        END
        AntennaGateArea 0.129 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.940 -0.210 3.080 0.210 ;
        RECT  2.680 -0.210 2.940 0.705 ;
        RECT  2.155 -0.210 2.680 0.210 ;
        RECT  1.985 -0.210 2.155 0.520 ;
        RECT  1.435 -0.210 1.985 0.210 ;
        RECT  1.265 -0.210 1.435 0.520 ;
        RECT  0.715 -0.210 1.265 0.210 ;
        RECT  0.545 -0.210 0.715 0.665 ;
        RECT  0.000 -0.210 0.545 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.815 2.310 3.080 2.730 ;
        RECT  2.645 2.060 2.815 2.730 ;
        RECT  0.825 2.310 2.645 2.730 ;
        RECT  0.655 1.800 0.825 2.730 ;
        RECT  0.000 2.310 0.655 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  1.520 0.900 1.780 1.200 ;
        RECT  0.600 0.900 1.520 1.020 ;
        RECT  0.480 0.785 0.600 1.635 ;
        RECT  0.355 0.785 0.480 0.905 ;
        RECT  0.455 1.515 0.480 1.635 ;
        RECT  0.285 1.515 0.455 1.945 ;
        RECT  0.185 0.435 0.355 0.905 ;
    END
END NOR3BX4AD
MACRO NOR3BXLAD
    CLASS CORE ;
    FOREIGN NOR3BXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.730 1.610 1.645 ;
        RECT  1.425 0.730 1.470 0.905 ;
        RECT  1.425 1.475 1.470 1.645 ;
        RECT  0.710 0.730 1.425 0.880 ;
        END
        AntennaDiffArea 0.19 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.000 0.770 1.420 ;
        END
        AntennaGateArea 0.0604 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.010 1.065 1.415 ;
        END
        AntennaGateArea 0.06 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.010 0.270 1.270 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.0424 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.185 -0.210 1.680 0.210 ;
        RECT  0.495 -0.210 1.185 0.325 ;
        RECT  0.000 -0.210 0.495 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.605 2.310 1.680 2.730 ;
        RECT  0.435 1.935 0.605 2.730 ;
        RECT  0.000 2.310 0.435 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.305 1.010 1.350 1.270 ;
        RECT  1.185 1.010 1.305 1.665 ;
        RECT  0.510 1.545 1.185 1.665 ;
        RECT  0.390 0.625 0.510 1.665 ;
        RECT  0.330 0.625 0.390 0.745 ;
        RECT  0.085 1.495 0.390 1.665 ;
        RECT  0.210 0.330 0.330 0.745 ;
        RECT  0.070 0.330 0.210 0.450 ;
    END
END NOR3BXLAD
MACRO NOR3X1AD
    CLASS CORE ;
    FOREIGN NOR3X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.690 1.330 1.740 ;
        RECT  1.190 0.690 1.230 1.955 ;
        RECT  0.095 0.690 1.190 0.860 ;
        RECT  1.060 1.525 1.190 1.955 ;
        END
        AntennaDiffArea 0.283 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 1.020 0.455 1.375 ;
        RECT  0.070 1.145 0.250 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.020 0.785 1.655 ;
        END
        AntennaGateArea 0.09 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.020 1.070 1.405 ;
        END
        AntennaGateArea 0.09 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 -0.210 1.400 0.210 ;
        RECT  1.055 -0.210 1.225 0.375 ;
        RECT  0.685 -0.210 1.055 0.210 ;
        RECT  0.515 -0.210 0.685 0.375 ;
        RECT  0.000 -0.210 0.515 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.305 2.310 1.400 2.730 ;
        RECT  0.135 1.495 0.305 2.730 ;
        RECT  0.000 2.310 0.135 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
	 END
END NOR3X1AD
MACRO NOR3X2AD
    CLASS CORE ;
    FOREIGN NOR3X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.195 0.415 1.365 2.055 ;
        RECT  1.190 0.745 1.195 2.055 ;
        RECT  0.645 0.745 1.190 0.905 ;
        RECT  1.075 1.625 1.190 2.055 ;
        RECT  0.475 0.415 0.645 0.905 ;
        END
        AntennaDiffArea 0.553 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.275 1.025 0.495 1.375 ;
        RECT  0.070 1.145 0.275 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.025 0.790 1.655 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.025 1.070 1.465 ;
        END
        AntennaGateArea 0.162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.005 -0.210 1.680 0.210 ;
        RECT  0.835 -0.210 1.005 0.625 ;
        RECT  0.285 -0.210 0.835 0.210 ;
        RECT  0.115 -0.210 0.285 0.845 ;
        RECT  0.000 -0.210 0.115 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.345 2.310 1.680 2.730 ;
        RECT  0.175 1.575 0.345 2.730 ;
        RECT  0.000 2.310 0.175 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
	 END
END NOR3X2AD
MACRO NOR3X4AD
    CLASS CORE ;
    FOREIGN NOR3X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.770 2.450 1.890 ;
        RECT  2.100 0.770 2.310 0.910 ;
        RECT  1.380 1.760 2.310 1.890 ;
        RECT  1.880 0.360 2.100 0.910 ;
        RECT  1.840 0.360 1.880 0.740 ;
        RECT  1.380 0.610 1.840 0.740 ;
        RECT  1.120 0.360 1.380 0.740 ;
        RECT  1.120 1.760 1.380 2.140 ;
        RECT  0.660 0.610 1.120 0.740 ;
        RECT  0.400 0.360 0.660 0.740 ;
        END
        AntennaDiffArea 0.782 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.030 2.150 1.640 ;
        RECT  0.490 1.520 2.030 1.640 ;
        RECT  0.350 1.010 0.490 1.640 ;
        RECT  0.320 1.010 0.350 1.270 ;
        END
        AntennaGateArea 0.324 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.020 1.820 1.280 ;
        RECT  1.620 0.860 1.740 1.280 ;
        RECT  1.095 0.860 1.620 0.980 ;
        RECT  0.740 0.860 1.095 1.050 ;
        RECT  0.620 0.860 0.740 1.270 ;
        END
        AntennaGateArea 0.324 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.215 1.100 1.475 1.330 ;
        RECT  1.145 1.170 1.215 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.415 -0.210 2.520 0.210 ;
        RECT  2.245 -0.210 2.415 0.650 ;
        RECT  1.695 -0.210 2.245 0.210 ;
        RECT  1.525 -0.210 1.695 0.490 ;
        RECT  0.975 -0.210 1.525 0.210 ;
        RECT  0.805 -0.210 0.975 0.490 ;
        RECT  0.255 -0.210 0.805 0.210 ;
        RECT  0.085 -0.210 0.255 0.780 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.340 2.310 2.520 2.730 ;
        RECT  2.080 2.010 2.340 2.730 ;
        RECT  0.230 2.310 2.080 2.730 ;
        RECT  0.090 1.570 0.230 2.730 ;
        RECT  0.000 2.310 0.090 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
	 END
END NOR3X4AD
MACRO NOR3X6AD
    CLASS CORE ;
    FOREIGN NOR3X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.740 0.410 3.815 0.840 ;
        RECT  3.600 0.410 3.740 1.925 ;
        RECT  1.460 0.410 3.600 0.540 ;
        RECT  3.475 1.450 3.600 1.925 ;
        RECT  2.825 1.750 3.475 1.925 ;
        RECT  1.405 1.775 2.825 1.925 ;
        RECT  1.290 0.410 1.460 0.705 ;
        RECT  1.235 1.775 1.405 1.990 ;
        RECT  0.485 0.575 1.290 0.705 ;
        END
        AntennaDiffArea 1.463 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.340 1.140 2.740 1.260 ;
        RECT  2.220 1.140 2.340 1.650 ;
        RECT  0.610 1.530 2.220 1.650 ;
        RECT  0.490 1.010 0.610 1.650 ;
        RECT  0.310 1.010 0.490 1.375 ;
        END
        AntennaGateArea 0.4828 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.035 0.900 3.155 1.280 ;
        RECT  1.970 0.900 3.035 1.020 ;
        RECT  1.850 0.900 1.970 1.410 ;
        RECT  1.690 1.125 1.850 1.410 ;
        RECT  0.890 1.290 1.690 1.410 ;
        RECT  0.760 1.020 0.890 1.410 ;
        END
        AntennaGateArea 0.4839 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.360 0.660 3.480 1.260 ;
        RECT  1.725 0.660 3.360 0.780 ;
        RECT  1.605 0.660 1.725 1.005 ;
        RECT  1.570 0.865 1.605 1.005 ;
        RECT  1.050 0.865 1.570 1.170 ;
        END
        AntennaGateArea 0.483 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.470 -0.210 3.920 0.210 ;
        RECT  3.210 -0.210 3.470 0.290 ;
        RECT  2.670 -0.210 3.210 0.210 ;
        RECT  2.410 -0.210 2.670 0.290 ;
        RECT  1.885 -0.210 2.410 0.210 ;
        RECT  1.625 -0.210 1.885 0.290 ;
        RECT  1.125 -0.210 1.625 0.210 ;
        RECT  0.865 -0.210 1.125 0.455 ;
        RECT  0.340 -0.210 0.865 0.210 ;
        RECT  0.170 -0.210 0.340 0.780 ;
        RECT  0.000 -0.210 0.170 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.585 2.310 3.920 2.730 ;
        RECT  2.415 2.045 2.585 2.730 ;
        RECT  0.370 2.310 2.415 2.730 ;
        RECT  0.200 1.495 0.370 2.730 ;
        RECT  0.000 2.310 0.200 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
	 END
END NOR3X6AD
MACRO NOR3X8AD
    CLASS CORE ;
    FOREIGN NOR3X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.900 1.005 5.110 1.515 ;
        RECT  4.650 0.670 4.900 2.085 ;
        RECT  4.375 0.670 4.650 0.880 ;
        RECT  1.170 1.825 4.650 2.085 ;
        RECT  4.205 0.420 4.375 0.880 ;
        RECT  3.655 0.670 4.205 0.880 ;
        RECT  3.485 0.410 3.655 0.880 ;
        RECT  0.615 0.410 3.485 0.550 ;
        RECT  0.445 0.410 0.615 0.850 ;
        END
        AntennaDiffArea 1.6 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.360 1.015 4.480 1.655 ;
        RECT  2.545 1.535 4.360 1.655 ;
        RECT  2.545 1.150 2.675 1.270 ;
        RECT  2.285 1.150 2.545 1.655 ;
        RECT  2.155 1.150 2.285 1.270 ;
        RECT  0.815 1.535 2.285 1.655 ;
        RECT  0.580 1.470 0.815 1.890 ;
        RECT  0.460 1.080 0.580 1.655 ;
        RECT  0.280 1.080 0.460 1.200 ;
        END
        AntennaGateArea 0.6428 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.995 1.010 4.115 1.410 ;
        RECT  3.040 1.290 3.995 1.410 ;
        RECT  2.920 0.910 3.040 1.410 ;
        RECT  1.985 0.910 2.920 1.030 ;
        RECT  1.750 0.910 1.985 1.410 ;
        RECT  1.055 1.290 1.750 1.410 ;
        RECT  0.935 1.150 1.055 1.410 ;
        RECT  0.820 1.150 0.935 1.270 ;
        RECT  0.700 1.010 0.820 1.270 ;
        END
        AntennaGateArea 0.6435 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.340 1.050 3.740 1.170 ;
        RECT  3.220 0.670 3.340 1.170 ;
        RECT  1.440 0.670 3.220 0.790 ;
        RECT  1.180 0.670 1.440 1.170 ;
        END
        AntennaGateArea 0.6435 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.735 -0.210 5.320 0.210 ;
        RECT  4.565 -0.210 4.735 0.550 ;
        RECT  4.015 -0.210 4.565 0.210 ;
        RECT  3.845 -0.210 4.015 0.550 ;
        RECT  3.320 -0.210 3.845 0.210 ;
        RECT  3.060 -0.210 3.320 0.290 ;
        RECT  2.560 -0.210 3.060 0.210 ;
        RECT  2.300 -0.210 2.560 0.290 ;
        RECT  1.800 -0.210 2.300 0.210 ;
        RECT  1.540 -0.210 1.800 0.290 ;
        RECT  1.040 -0.210 1.540 0.210 ;
        RECT  0.780 -0.210 1.040 0.290 ;
        RECT  0.255 -0.210 0.780 0.210 ;
        RECT  0.085 -0.210 0.255 0.850 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.725 2.310 5.320 2.730 ;
        RECT  4.555 2.205 4.725 2.730 ;
        RECT  2.495 2.310 4.555 2.730 ;
        RECT  2.325 2.205 2.495 2.730 ;
        RECT  0.340 2.310 2.325 2.730 ;
        RECT  0.195 1.375 0.340 2.730 ;
        RECT  0.000 2.310 0.195 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.320 2.520 ;
	 END
END NOR3X8AD
MACRO NOR3XLAD
    CLASS CORE ;
    FOREIGN NOR3XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.735 1.330 1.695 ;
        RECT  0.095 0.735 1.190 0.905 ;
        RECT  1.060 1.525 1.190 1.695 ;
        END
        AntennaDiffArea 0.19 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 1.025 0.455 1.375 ;
        RECT  0.070 1.145 0.250 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.025 0.785 1.655 ;
        END
        AntennaGateArea 0.06 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.025 1.070 1.405 ;
        END
        AntennaGateArea 0.0604 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.225 -0.210 1.400 0.210 ;
        RECT  1.055 -0.210 1.225 0.375 ;
        RECT  0.685 -0.210 1.055 0.210 ;
        RECT  0.515 -0.210 0.685 0.375 ;
        RECT  0.000 -0.210 0.515 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.305 2.310 1.400 2.730 ;
        RECT  0.135 1.495 0.305 2.730 ;
        RECT  0.000 2.310 0.135 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
	 END
END NOR3XLAD
MACRO NOR4BBX1AD
    CLASS CORE ;
    FOREIGN NOR4BBX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.640 2.730 1.690 ;
        RECT  1.580 0.640 2.590 0.780 ;
        RECT  2.575 1.550 2.590 1.690 ;
        RECT  2.435 1.550 2.575 2.070 ;
        RECT  1.460 0.640 1.580 0.900 ;
        END
        AntennaDiffArea 0.292 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.865 1.340 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.020 1.770 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.995 0.805 1.375 ;
        END
        AntennaGateArea 0.0474 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.015 0.250 1.275 ;
        RECT  0.070 1.015 0.210 1.375 ;
        END
        AntennaGateArea 0.0474 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.660 -0.210 2.800 0.210 ;
        RECT  1.800 -0.210 2.660 0.330 ;
        RECT  1.110 -0.210 1.800 0.210 ;
        RECT  0.550 -0.210 1.110 0.330 ;
        RECT  0.000 -0.210 0.550 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 2.310 2.800 2.730 ;
        RECT  1.070 1.975 1.370 2.095 ;
        RECT  0.810 1.975 1.070 2.730 ;
        RECT  0.510 1.975 0.810 2.095 ;
        RECT  0.000 2.310 0.810 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.310 1.020 2.415 1.280 ;
        RECT  2.190 1.020 2.310 1.855 ;
        RECT  0.490 1.735 2.190 1.855 ;
        RECT  1.950 1.020 2.070 1.615 ;
        RECT  1.055 1.495 1.950 1.615 ;
        RECT  0.935 0.750 1.055 1.615 ;
        RECT  0.730 0.750 0.935 0.870 ;
        RECT  0.840 1.495 0.935 1.615 ;
        RECT  0.370 0.725 0.490 1.855 ;
        RECT  0.095 0.725 0.370 0.895 ;
        RECT  0.080 1.495 0.370 1.675 ;
    END
END NOR4BBX1AD
MACRO NOR4BBX2AD
    CLASS CORE ;
    FOREIGN NOR4BBX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.460 1.980 1.630 2.150 ;
        RECT  0.220 1.980 1.460 2.100 ;
        RECT  1.245 0.330 1.365 0.850 ;
        RECT  0.710 0.625 1.245 0.745 ;
        RECT  0.450 0.335 0.710 0.745 ;
        RECT  0.190 0.625 0.450 0.745 ;
        RECT  0.190 1.425 0.220 2.100 ;
        RECT  0.070 0.625 0.190 2.100 ;
        END
        AntennaDiffArea 0.604 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.605 1.040 2.665 1.300 ;
        RECT  2.485 1.040 2.605 1.860 ;
        RECT  0.490 1.740 2.485 1.860 ;
        RECT  0.370 0.865 0.490 1.860 ;
        RECT  0.340 0.865 0.370 1.095 ;
        END
        AntennaGateArea 0.255 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 1.040 2.365 1.620 ;
        RECT  1.985 1.470 2.245 1.620 ;
        RECT  0.795 1.500 1.985 1.620 ;
        RECT  0.675 1.010 0.795 1.620 ;
        END
        AntennaGateArea 0.255 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.025 0.865 3.290 1.270 ;
        END
        AntennaGateArea 0.1074 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.410 0.865 3.580 1.335 ;
        END
        AntennaGateArea 0.112 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.205 -0.210 3.920 0.210 ;
        RECT  3.035 -0.210 3.205 0.400 ;
        RECT  1.795 -0.210 3.035 0.210 ;
        RECT  1.535 -0.210 1.795 0.400 ;
        RECT  1.030 -0.210 1.535 0.210 ;
        RECT  0.860 -0.210 1.030 0.505 ;
        RECT  0.305 -0.210 0.860 0.210 ;
        RECT  0.135 -0.210 0.305 0.505 ;
        RECT  0.000 -0.210 0.135 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.520 2.310 3.920 2.730 ;
        RECT  3.400 1.475 3.520 2.730 ;
        RECT  3.260 1.475 3.400 1.595 ;
        RECT  2.955 2.310 3.400 2.730 ;
        RECT  2.695 2.230 2.955 2.730 ;
        RECT  0.340 2.310 2.695 2.730 ;
        RECT  0.080 2.220 0.340 2.730 ;
        RECT  0.000 2.310 0.080 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  3.730 0.520 3.850 2.010 ;
        RECT  1.630 0.520 3.730 0.640 ;
        RECT  3.690 1.430 3.730 2.010 ;
        RECT  3.140 1.775 3.205 1.945 ;
        RECT  3.020 1.595 3.140 1.945 ;
        RECT  2.905 1.595 3.020 1.715 ;
        RECT  2.785 0.760 2.905 1.715 ;
        RECT  2.065 0.760 2.785 0.880 ;
        RECT  1.945 0.760 2.065 1.300 ;
        RECT  1.870 1.180 1.945 1.300 ;
        RECT  1.750 1.180 1.870 1.380 ;
        RECT  1.155 1.260 1.750 1.380 ;
        RECT  1.510 0.520 1.630 1.140 ;
        RECT  1.370 1.020 1.510 1.140 ;
        RECT  1.035 1.010 1.155 1.380 ;
    END
END NOR4BBX2AD
MACRO NOR4BBX4AD
    CLASS CORE ;
    FOREIGN NOR4BBX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.300 0.640 3.440 1.695 ;
        RECT  0.740 0.640 3.300 0.780 ;
        RECT  3.010 1.555 3.300 1.695 ;
        RECT  2.870 1.555 3.010 2.075 ;
        RECT  2.060 1.760 2.870 1.900 ;
        RECT  1.800 1.760 2.060 2.175 ;
        END
        AntennaDiffArea 0.817 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.060 1.020 3.180 1.430 ;
        RECT  2.720 1.310 3.060 1.430 ;
        RECT  2.600 1.310 2.720 1.640 ;
        RECT  0.860 1.520 2.600 1.640 ;
        RECT  0.585 1.140 0.860 1.640 ;
        END
        AntennaGateArea 0.27 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.070 2.900 1.190 ;
        RECT  2.320 1.070 2.440 1.400 ;
        RECT  1.330 1.280 2.320 1.400 ;
        RECT  1.190 1.140 1.330 1.400 ;
        RECT  0.980 1.140 1.190 1.260 ;
        END
        AntennaGateArea 0.2709 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.710 1.705 3.850 2.190 ;
        RECT  3.450 2.070 3.710 2.190 ;
        END
        AntennaGateArea 0.1304 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.160 0.330 0.535 0.535 ;
        END
        AntennaGateArea 0.128 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.260 -0.210 3.920 0.210 ;
        RECT  2.740 -0.210 3.260 0.230 ;
        RECT  2.020 -0.210 2.740 0.210 ;
        RECT  1.760 -0.210 2.020 0.230 ;
        RECT  1.195 -0.210 1.760 0.210 ;
        RECT  0.675 -0.210 1.195 0.230 ;
        RECT  0.000 -0.210 0.675 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.330 2.310 3.920 2.730 ;
        RECT  3.210 1.820 3.330 2.730 ;
        RECT  0.695 2.310 3.210 2.730 ;
        RECT  0.525 1.760 0.695 2.730 ;
        RECT  0.000 2.310 0.525 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  3.690 0.380 3.810 1.585 ;
        RECT  2.590 0.380 3.690 0.500 ;
        RECT  3.565 1.415 3.690 1.585 ;
        RECT  2.330 0.330 2.590 0.500 ;
        RECT  1.570 0.380 2.330 0.500 ;
        RECT  1.825 1.040 2.185 1.160 ;
        RECT  1.625 0.900 1.825 1.160 ;
        RECT  0.310 0.900 1.625 1.020 ;
        RECT  1.310 0.330 1.570 0.500 ;
        RECT  0.175 0.700 0.310 2.175 ;
        RECT  0.085 0.700 0.175 0.870 ;
    END
END NOR4BBX4AD
MACRO NOR4BBXLAD
    CLASS CORE ;
    FOREIGN NOR4BBXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.730 2.730 1.810 ;
        RECT  1.580 0.730 2.590 0.870 ;
        RECT  2.430 1.550 2.590 1.810 ;
        RECT  1.460 0.680 1.580 0.940 ;
        END
        AntennaDiffArea 0.205 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.865 1.340 1.375 ;
        END
        AntennaGateArea 0.0644 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.060 1.770 1.375 ;
        END
        AntennaGateArea 0.064 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.995 0.805 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.015 0.250 1.275 ;
        RECT  0.070 1.015 0.210 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.660 -0.210 2.800 0.210 ;
        RECT  1.800 -0.210 2.660 0.330 ;
        RECT  1.110 -0.210 1.800 0.210 ;
        RECT  0.550 -0.210 1.110 0.330 ;
        RECT  0.000 -0.210 0.550 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.070 2.310 2.800 2.730 ;
        RECT  1.070 1.975 1.365 2.095 ;
        RECT  0.810 1.975 1.070 2.730 ;
        RECT  0.505 1.975 0.810 2.095 ;
        RECT  0.000 2.310 0.810 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.310 1.020 2.415 1.280 ;
        RECT  2.190 1.020 2.310 1.855 ;
        RECT  0.490 1.735 2.190 1.855 ;
        RECT  1.950 1.020 2.070 1.615 ;
        RECT  1.055 1.495 1.950 1.615 ;
        RECT  0.935 0.750 1.055 1.615 ;
        RECT  0.730 0.750 0.935 0.870 ;
        RECT  0.840 1.495 0.935 1.615 ;
        RECT  0.370 0.725 0.490 1.855 ;
        RECT  0.095 0.725 0.370 0.895 ;
        RECT  0.080 1.495 0.370 1.675 ;
    END
END NOR4BBXLAD
MACRO NOR4BX1AD
    CLASS CORE ;
    FOREIGN NOR4BX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.575 2.170 1.905 ;
        RECT  0.980 0.575 2.030 0.745 ;
        RECT  1.790 1.735 2.030 1.905 ;
        RECT  0.810 0.575 0.980 0.810 ;
        END
        AntennaDiffArea 0.3 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.000 0.785 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.010 1.185 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.865 1.610 1.270 ;
        END
        AntennaGateArea 0.09 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.995 0.490 1.375 ;
        END
        AntennaGateArea 0.0472 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.010 -0.210 2.240 0.210 ;
        RECT  1.230 -0.210 2.010 0.315 ;
        RECT  0.620 -0.210 1.230 0.210 ;
        RECT  0.450 -0.210 0.620 0.860 ;
        RECT  0.000 -0.210 0.450 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.715 2.310 2.240 2.730 ;
        RECT  0.545 1.735 0.715 2.730 ;
        RECT  0.000 2.310 0.545 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.735 1.010 1.855 1.615 ;
        RECT  0.190 1.495 1.735 1.615 ;
        RECT  0.190 0.690 0.260 0.860 ;
        RECT  0.070 0.690 0.190 1.615 ;
    END
END NOR4BX1AD
MACRO NOR4BX2AD
    CLASS CORE ;
    FOREIGN NOR4BX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.460 1.980 1.630 2.150 ;
        RECT  0.220 1.980 1.460 2.100 ;
        RECT  0.190 0.550 1.435 0.670 ;
        RECT  0.190 1.425 0.220 2.100 ;
        RECT  0.070 0.550 0.190 2.100 ;
        END
        AntennaDiffArea 0.604 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.605 1.025 2.665 1.285 ;
        RECT  2.485 1.025 2.605 1.860 ;
        RECT  0.490 1.740 2.485 1.860 ;
        RECT  0.370 0.865 0.490 1.860 ;
        RECT  0.340 0.865 0.370 1.095 ;
        END
        AntennaGateArea 0.255 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.245 1.040 2.365 1.620 ;
        RECT  1.985 1.470 2.245 1.620 ;
        RECT  0.795 1.500 1.985 1.620 ;
        RECT  0.675 1.030 0.795 1.620 ;
        END
        AntennaGateArea 0.255 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.040 2.065 1.300 ;
        RECT  1.750 1.040 1.890 1.380 ;
        RECT  1.155 1.260 1.750 1.380 ;
        RECT  1.035 1.030 1.155 1.380 ;
        END
        AntennaGateArea 0.255 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.820 1.025 3.050 1.375 ;
        END
        AntennaGateArea 0.1124 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.915 -0.210 3.360 0.210 ;
        RECT  2.745 -0.210 2.915 0.665 ;
        RECT  1.795 -0.210 2.745 0.210 ;
        RECT  1.535 -0.210 1.795 0.390 ;
        RECT  1.030 -0.210 1.535 0.210 ;
        RECT  0.860 -0.210 1.030 0.430 ;
        RECT  0.305 -0.210 0.860 0.210 ;
        RECT  0.135 -0.210 0.305 0.430 ;
        RECT  0.000 -0.210 0.135 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.845 2.310 3.360 2.730 ;
        RECT  2.725 1.525 2.845 2.730 ;
        RECT  0.340 2.310 2.725 2.730 ;
        RECT  0.080 2.220 0.340 2.730 ;
        RECT  0.000 2.310 0.080 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  3.250 0.495 3.290 1.735 ;
        RECT  3.170 0.495 3.250 1.985 ;
        RECT  3.105 0.495 3.170 0.665 ;
        RECT  1.630 0.785 3.170 0.905 ;
        RECT  3.080 1.495 3.170 1.985 ;
        RECT  1.510 0.785 1.630 1.140 ;
        RECT  1.370 1.020 1.510 1.140 ;
    END
END NOR4BX2AD
MACRO NOR4BX4AD
    CLASS CORE ;
    FOREIGN NOR4BX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.160 0.560 3.290 1.985 ;
        RECT  2.685 0.560 3.160 0.770 ;
        RECT  2.925 1.865 3.160 1.985 ;
        RECT  2.805 1.865 2.925 2.140 ;
        RECT  1.720 2.020 2.805 2.140 ;
        RECT  0.710 0.560 2.685 0.680 ;
        END
        AntennaDiffArea 0.803 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.920 1.010 3.040 1.745 ;
        RECT  2.685 1.625 2.920 1.745 ;
        RECT  2.565 1.625 2.685 1.900 ;
        RECT  0.785 1.780 2.565 1.900 ;
        RECT  0.615 1.085 0.785 1.900 ;
        END
        AntennaGateArea 0.27 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.620 1.000 2.740 1.505 ;
        RECT  2.445 1.385 2.620 1.505 ;
        RECT  2.325 1.385 2.445 1.660 ;
        RECT  1.145 1.540 2.325 1.660 ;
        RECT  1.025 1.085 1.145 1.660 ;
        RECT  0.910 1.085 1.025 1.375 ;
        END
        AntennaGateArea 0.2709 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.430 1.265 ;
        RECT  2.170 1.145 2.310 1.265 ;
        RECT  2.030 1.145 2.170 1.420 ;
        RECT  1.450 1.300 2.030 1.420 ;
        RECT  1.330 1.040 1.450 1.420 ;
        END
        AntennaGateArea 0.3209 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.975 0.230 1.375 ;
        END
        AntennaGateArea 0.16 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.110 -0.210 3.360 0.210 ;
        RECT  2.640 -0.210 3.110 0.255 ;
        RECT  2.015 -0.210 2.640 0.210 ;
        RECT  1.845 -0.210 2.015 0.255 ;
        RECT  1.095 -0.210 1.845 0.210 ;
        RECT  0.625 -0.210 1.095 0.255 ;
        RECT  0.000 -0.210 0.625 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.215 2.310 3.360 2.730 ;
        RECT  3.045 2.105 3.215 2.730 ;
        RECT  0.655 2.310 3.045 2.730 ;
        RECT  0.485 2.035 0.655 2.730 ;
        RECT  0.000 2.310 0.485 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  1.650 0.800 1.910 1.180 ;
        RECT  0.470 0.800 1.650 0.920 ;
        RECT  0.350 0.670 0.470 1.615 ;
        RECT  0.255 0.670 0.350 0.790 ;
        RECT  0.275 1.495 0.350 1.615 ;
        RECT  0.105 1.495 0.275 2.185 ;
        RECT  0.085 0.360 0.255 0.790 ;
    END
END NOR4BX4AD
MACRO NOR4BXLAD
    CLASS CORE ;
    FOREIGN NOR4BXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.705 2.170 1.875 ;
        RECT  0.765 0.705 2.030 0.845 ;
        RECT  1.745 1.735 2.030 1.875 ;
        END
        AntennaDiffArea 0.209 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.000 0.785 1.375 ;
        END
        AntennaGateArea 0.064 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.010 1.185 1.375 ;
        END
        AntennaGateArea 0.064 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.990 1.610 1.375 ;
        END
        AntennaGateArea 0.064 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.995 0.490 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.010 -0.210 2.240 0.210 ;
        RECT  1.230 -0.210 2.010 0.315 ;
        RECT  0.620 -0.210 1.230 0.210 ;
        RECT  0.450 -0.210 0.620 0.860 ;
        RECT  0.000 -0.210 0.450 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.760 2.310 2.240 2.730 ;
        RECT  0.500 1.735 0.760 2.730 ;
        RECT  0.000 2.310 0.500 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.735 1.010 1.855 1.615 ;
        RECT  0.190 1.495 1.735 1.615 ;
        RECT  0.190 0.690 0.260 0.860 ;
        RECT  0.070 0.690 0.190 1.615 ;
    END
END NOR4BXLAD
MACRO NOR4X1AD
    CLASS CORE ;
    FOREIGN NOR4X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.355 1.425 1.525 1.980 ;
        RECT  1.290 1.425 1.355 1.655 ;
        RECT  1.170 0.655 1.290 1.655 ;
        RECT  1.115 0.655 1.170 0.995 ;
        RECT  0.565 0.875 1.115 0.995 ;
        RECT  0.395 0.655 0.565 0.995 ;
        END
        AntennaDiffArea 0.292 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.590 0.230 1.285 ;
        END
        AntennaGateArea 0.09 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.115 0.760 1.375 ;
        END
        AntennaGateArea 0.0906 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.115 1.050 1.650 ;
        END
        AntennaGateArea 0.0906 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.465 0.605 1.610 1.285 ;
        END
        AntennaGateArea 0.09 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 -0.210 1.680 0.210 ;
        RECT  1.345 -0.210 1.515 0.350 ;
        RECT  0.970 -0.210 1.345 0.210 ;
        RECT  0.710 -0.210 0.970 0.755 ;
        RECT  0.335 -0.210 0.710 0.210 ;
        RECT  0.165 -0.210 0.335 0.350 ;
        RECT  0.000 -0.210 0.165 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.325 2.310 1.680 2.730 ;
        RECT  0.155 1.495 0.325 2.730 ;
        RECT  0.000 2.310 0.155 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
	 END
END NOR4X1AD
MACRO NOR4X2AD
    CLASS CORE ;
    FOREIGN NOR4X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.410 1.930 1.580 2.100 ;
        RECT  0.575 1.930 1.410 2.050 ;
        RECT  0.190 0.550 1.385 0.670 ;
        RECT  0.455 1.890 0.575 2.050 ;
        RECT  0.210 1.890 0.455 2.010 ;
        RECT  0.190 1.425 0.210 2.010 ;
        RECT  0.070 0.550 0.190 2.010 ;
        END
        AntennaDiffArea 0.604 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.510 0.510 2.630 1.285 ;
        RECT  1.625 0.510 2.510 0.630 ;
        RECT  1.505 0.510 1.625 0.910 ;
        RECT  0.490 0.790 1.505 0.910 ;
        RECT  0.320 0.790 0.490 1.270 ;
        END
        AntennaGateArea 0.255 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.230 0.765 2.390 0.885 ;
        RECT  2.110 0.765 2.230 1.810 ;
        RECT  2.030 1.425 2.110 1.810 ;
        RECT  0.790 1.690 2.030 1.810 ;
        RECT  0.670 1.030 0.790 1.810 ;
        RECT  0.625 1.030 0.670 1.290 ;
        END
        AntennaGateArea 0.255 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 0.785 1.910 1.570 ;
        RECT  1.050 1.450 1.790 1.570 ;
        RECT  1.050 1.030 1.105 1.290 ;
        RECT  0.910 1.030 1.050 1.570 ;
        END
        AntennaGateArea 0.255 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.030 1.655 1.330 ;
        END
        AntennaGateArea 0.255 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.745 -0.210 2.800 0.210 ;
        RECT  1.485 -0.210 1.745 0.390 ;
        RECT  0.980 -0.210 1.485 0.210 ;
        RECT  0.810 -0.210 0.980 0.430 ;
        RECT  0.255 -0.210 0.810 0.210 ;
        RECT  0.085 -0.210 0.255 0.430 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.715 2.310 2.800 2.730 ;
        RECT  2.545 1.420 2.715 2.730 ;
        RECT  0.360 2.310 2.545 2.730 ;
        RECT  0.100 2.130 0.360 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
	 END
END NOR4X2AD
MACRO NOR4X4AD
    CLASS CORE ;
    FOREIGN NOR4X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.295 0.560 5.415 2.010 ;
        RECT  4.305 0.560 5.295 0.680 ;
        RECT  5.055 1.890 5.295 2.010 ;
        RECT  4.935 1.890 5.055 2.050 ;
        RECT  4.035 1.930 4.935 2.050 ;
        RECT  4.185 0.330 4.305 0.680 ;
        RECT  3.525 1.930 4.035 2.170 ;
        RECT  3.070 1.930 3.525 2.050 ;
        RECT  2.950 1.450 3.070 2.050 ;
        RECT  2.525 1.450 2.950 1.570 ;
        RECT  2.405 1.450 2.525 2.050 ;
        RECT  1.575 1.930 2.405 2.050 ;
        RECT  1.405 1.930 1.575 2.100 ;
        RECT  0.570 1.930 1.405 2.050 ;
        RECT  1.190 0.410 1.310 0.670 ;
        RECT  0.190 0.550 1.190 0.670 ;
        RECT  0.450 1.890 0.570 2.050 ;
        RECT  0.190 1.890 0.450 2.010 ;
        RECT  0.070 0.550 0.190 2.010 ;
        END
        AntennaDiffArea 1.199 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.055 0.800 5.175 1.270 ;
        RECT  4.060 0.800 5.055 0.920 ;
        RECT  3.940 0.410 4.060 0.920 ;
        RECT  1.550 0.410 3.940 0.530 ;
        RECT  1.430 0.410 1.550 0.910 ;
        RECT  0.490 0.790 1.430 0.910 ;
        RECT  0.320 0.790 0.490 1.270 ;
        END
        AntennaGateArea 0.503 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.695 1.040 4.815 1.720 ;
        RECT  3.340 1.600 4.695 1.720 ;
        RECT  3.220 1.190 3.340 1.720 ;
        RECT  2.495 1.190 3.220 1.310 ;
        RECT  2.270 1.130 2.495 1.330 ;
        RECT  2.150 1.130 2.270 1.810 ;
        RECT  0.790 1.690 2.150 1.810 ;
        RECT  0.670 1.030 0.790 1.810 ;
        RECT  0.620 1.030 0.670 1.290 ;
        END
        AntennaGateArea 0.5043 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.385 1.040 4.505 1.480 ;
        RECT  3.580 1.360 4.385 1.480 ;
        RECT  3.460 0.890 3.580 1.480 ;
        RECT  2.030 0.890 3.460 1.010 ;
        RECT  1.910 0.890 2.030 1.570 ;
        RECT  1.050 1.450 1.910 1.570 ;
        RECT  1.050 1.030 1.100 1.290 ;
        RECT  0.910 1.030 1.050 1.570 ;
        END
        AntennaGateArea 0.505 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.820 1.100 3.995 1.220 ;
        RECT  3.700 0.650 3.820 1.220 ;
        RECT  1.790 0.650 3.700 0.770 ;
        RECT  1.670 0.650 1.790 1.330 ;
        RECT  1.360 1.110 1.670 1.330 ;
        END
        AntennaGateArea 0.505 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.410 -0.210 5.600 0.210 ;
        RECT  5.240 -0.210 5.410 0.430 ;
        RECT  4.690 -0.210 5.240 0.210 ;
        RECT  4.520 -0.210 4.690 0.415 ;
        RECT  3.945 -0.210 4.520 0.210 ;
        RECT  3.685 -0.210 3.945 0.290 ;
        RECT  1.810 -0.210 3.685 0.210 ;
        RECT  1.550 -0.210 1.810 0.290 ;
        RECT  0.975 -0.210 1.550 0.210 ;
        RECT  0.805 -0.210 0.975 0.430 ;
        RECT  0.255 -0.210 0.805 0.210 ;
        RECT  0.085 -0.210 0.255 0.430 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.435 2.310 5.600 2.730 ;
        RECT  5.175 2.130 5.435 2.730 ;
        RECT  2.815 2.310 5.175 2.730 ;
        RECT  2.645 1.690 2.815 2.730 ;
        RECT  0.360 2.310 2.645 2.730 ;
        RECT  0.100 2.130 0.360 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
	 END
END NOR4X4AD
MACRO NOR4X6AD
    CLASS CORE ;
    FOREIGN NOR4X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.005 0.535 8.075 1.380 ;
        RECT  7.860 0.535 8.005 2.120 ;
        RECT  7.645 0.535 7.860 0.715 ;
        RECT  7.835 1.170 7.860 2.120 ;
        RECT  7.285 1.170 7.835 1.380 ;
        RECT  7.475 0.345 7.645 0.715 ;
        RECT  6.925 0.535 7.475 0.715 ;
        RECT  7.115 1.170 7.285 1.860 ;
        RECT  6.565 1.170 7.115 1.380 ;
        RECT  6.755 0.345 6.925 0.715 ;
        RECT  6.205 0.535 6.755 0.715 ;
        RECT  6.395 1.170 6.565 1.860 ;
        RECT  6.035 0.345 6.205 0.715 ;
        RECT  5.485 0.535 6.035 0.715 ;
        RECT  5.315 0.345 5.485 0.715 ;
        RECT  4.765 0.535 5.315 0.715 ;
        RECT  4.595 0.345 4.765 0.715 ;
        RECT  4.045 0.535 4.595 0.715 ;
        RECT  3.875 0.345 4.045 0.715 ;
        RECT  3.325 0.535 3.875 0.715 ;
        RECT  3.155 0.345 3.325 0.715 ;
        RECT  2.605 0.535 3.155 0.715 ;
        RECT  2.435 0.345 2.605 0.715 ;
        RECT  1.885 0.535 2.435 0.715 ;
        RECT  1.715 0.345 1.885 0.715 ;
        RECT  1.165 0.535 1.715 0.715 ;
        RECT  0.995 0.345 1.165 0.715 ;
        END
        AntennaDiffArea 1.966 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.385 0.845 2.345 0.965 ;
        RECT  0.865 0.845 1.385 1.050 ;
        END
        AntennaGateArea 0.81 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.665 0.840 4.185 1.050 ;
        RECT  2.670 0.840 3.665 0.960 ;
        END
        AntennaGateArea 0.81 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.295 0.840 5.960 0.960 ;
        RECT  4.785 0.840 5.295 1.050 ;
        RECT  4.500 0.840 4.785 0.960 ;
        END
        AntennaGateArea 0.81 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.695 0.840 7.740 0.960 ;
        RECT  6.185 0.840 6.695 1.050 ;
        END
        AntennaGateArea 0.81 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.005 -0.210 8.680 0.210 ;
        RECT  7.835 -0.210 8.005 0.415 ;
        RECT  7.285 -0.210 7.835 0.210 ;
        RECT  7.115 -0.210 7.285 0.415 ;
        RECT  6.565 -0.210 7.115 0.210 ;
        RECT  6.395 -0.210 6.565 0.415 ;
        RECT  5.845 -0.210 6.395 0.210 ;
        RECT  5.675 -0.210 5.845 0.415 ;
        RECT  5.125 -0.210 5.675 0.210 ;
        RECT  4.955 -0.210 5.125 0.415 ;
        RECT  4.405 -0.210 4.955 0.210 ;
        RECT  4.235 -0.210 4.405 0.415 ;
        RECT  3.685 -0.210 4.235 0.210 ;
        RECT  3.515 -0.210 3.685 0.415 ;
        RECT  2.965 -0.210 3.515 0.210 ;
        RECT  2.795 -0.210 2.965 0.415 ;
        RECT  2.245 -0.210 2.795 0.210 ;
        RECT  2.075 -0.210 2.245 0.415 ;
        RECT  1.525 -0.210 2.075 0.210 ;
        RECT  1.355 -0.210 1.525 0.415 ;
        RECT  0.805 -0.210 1.355 0.210 ;
        RECT  0.635 -0.210 0.805 0.415 ;
        RECT  0.000 -0.210 0.635 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.245 2.310 8.680 2.730 ;
        RECT  2.075 1.585 2.245 2.730 ;
        RECT  1.525 2.310 2.075 2.730 ;
        RECT  1.355 1.585 1.525 2.730 ;
        RECT  0.805 2.310 1.355 2.730 ;
        RECT  0.635 1.325 0.805 2.730 ;
        RECT  0.000 2.310 0.635 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.680 2.520 ;
        LAYER M1 ;
        RECT  7.475 1.500 7.645 2.190 ;
        RECT  6.925 2.000 7.475 2.140 ;
        RECT  6.755 1.500 6.925 2.190 ;
        RECT  6.205 2.000 6.755 2.140 ;
        RECT  6.035 1.170 6.205 2.140 ;
        RECT  5.485 1.170 6.035 1.310 ;
        RECT  5.675 1.450 5.845 2.140 ;
        RECT  5.125 2.000 5.675 2.140 ;
        RECT  5.315 1.170 5.485 1.860 ;
        RECT  4.765 1.170 5.315 1.310 ;
        RECT  4.955 1.450 5.125 2.140 ;
        RECT  4.405 2.000 4.955 2.140 ;
        RECT  4.595 1.170 4.765 1.860 ;
        RECT  4.235 1.170 4.405 2.140 ;
        RECT  3.685 1.170 4.235 1.310 ;
        RECT  3.875 1.450 4.045 2.140 ;
        RECT  3.325 2.000 3.875 2.140 ;
        RECT  3.515 1.170 3.685 1.860 ;
        RECT  2.965 1.170 3.515 1.310 ;
        RECT  3.155 1.450 3.325 2.140 ;
        RECT  2.605 2.000 3.155 2.140 ;
        RECT  2.795 1.170 2.965 1.860 ;
        RECT  2.435 1.170 2.605 2.140 ;
        RECT  1.885 1.170 2.435 1.310 ;
        RECT  1.715 1.170 1.885 1.995 ;
        RECT  1.165 1.170 1.715 1.310 ;
        RECT  0.995 1.170 1.165 1.995 ;
    END
END NOR4X6AD
MACRO NOR4X8AD
    CLASS CORE ;
    FOREIGN NOR4X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.885 0.535 11.035 1.470 ;
        RECT  10.715 0.535 10.885 2.060 ;
        RECT  10.690 0.535 10.715 1.470 ;
        RECT  10.525 0.535 10.690 0.715 ;
        RECT  10.525 1.050 10.690 1.470 ;
        RECT  10.355 0.345 10.525 0.715 ;
        RECT  10.165 1.170 10.525 1.470 ;
        RECT  9.805 0.535 10.355 0.715 ;
        RECT  9.995 1.170 10.165 1.860 ;
        RECT  9.445 1.170 9.995 1.415 ;
        RECT  9.635 0.345 9.805 0.715 ;
        RECT  9.085 0.535 9.635 0.715 ;
        RECT  9.275 1.170 9.445 1.860 ;
        RECT  8.725 1.170 9.275 1.415 ;
        RECT  8.915 0.345 9.085 0.715 ;
        RECT  8.365 0.535 8.915 0.715 ;
        RECT  8.555 1.170 8.725 1.860 ;
        RECT  8.195 0.345 8.365 0.715 ;
        RECT  7.645 0.535 8.195 0.715 ;
        RECT  7.475 0.345 7.645 0.715 ;
        RECT  6.925 0.535 7.475 0.715 ;
        RECT  6.755 0.345 6.925 0.715 ;
        RECT  6.205 0.535 6.755 0.715 ;
        RECT  6.035 0.345 6.205 0.715 ;
        RECT  5.485 0.535 6.035 0.715 ;
        RECT  5.315 0.345 5.485 0.715 ;
        RECT  4.765 0.535 5.315 0.715 ;
        RECT  4.595 0.345 4.765 0.715 ;
        RECT  4.045 0.535 4.595 0.715 ;
        RECT  3.875 0.345 4.045 0.715 ;
        RECT  3.325 0.535 3.875 0.715 ;
        RECT  3.155 0.345 3.325 0.715 ;
        RECT  2.605 0.535 3.155 0.715 ;
        RECT  2.435 0.345 2.605 0.715 ;
        RECT  1.885 0.535 2.435 0.715 ;
        RECT  1.715 0.345 1.885 0.715 ;
        RECT  1.165 0.535 1.715 0.715 ;
        RECT  0.995 0.345 1.165 0.715 ;
        END
        AntennaDiffArea 2.649 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.935 0.840 3.080 0.960 ;
        RECT  1.425 0.840 1.935 1.050 ;
        RECT  1.020 0.840 1.425 0.960 ;
        END
        AntennaGateArea 1.12 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.735 0.840 5.460 0.960 ;
        RECT  4.225 0.840 4.735 1.050 ;
        RECT  3.400 0.840 4.225 0.960 ;
        END
        AntennaGateArea 1.12 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.255 0.840 8.120 0.960 ;
        RECT  6.745 0.840 7.255 1.050 ;
        RECT  6.060 0.840 6.745 0.960 ;
        END
        AntennaGateArea 1.12 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.935 0.840 10.385 0.960 ;
        RECT  8.425 0.840 8.935 1.050 ;
        END
        AntennaGateArea 1.12 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.885 -0.210 11.480 0.210 ;
        RECT  10.715 -0.210 10.885 0.415 ;
        RECT  10.165 -0.210 10.715 0.210 ;
        RECT  9.995 -0.210 10.165 0.415 ;
        RECT  9.445 -0.210 9.995 0.210 ;
        RECT  9.275 -0.210 9.445 0.415 ;
        RECT  8.725 -0.210 9.275 0.210 ;
        RECT  8.555 -0.210 8.725 0.415 ;
        RECT  8.005 -0.210 8.555 0.210 ;
        RECT  7.835 -0.210 8.005 0.415 ;
        RECT  7.285 -0.210 7.835 0.210 ;
        RECT  7.115 -0.210 7.285 0.415 ;
        RECT  6.565 -0.210 7.115 0.210 ;
        RECT  6.395 -0.210 6.565 0.415 ;
        RECT  5.845 -0.210 6.395 0.210 ;
        RECT  5.675 -0.210 5.845 0.415 ;
        RECT  5.125 -0.210 5.675 0.210 ;
        RECT  4.955 -0.210 5.125 0.415 ;
        RECT  4.405 -0.210 4.955 0.210 ;
        RECT  4.235 -0.210 4.405 0.415 ;
        RECT  3.685 -0.210 4.235 0.210 ;
        RECT  3.515 -0.210 3.685 0.415 ;
        RECT  2.965 -0.210 3.515 0.210 ;
        RECT  2.795 -0.210 2.965 0.415 ;
        RECT  2.245 -0.210 2.795 0.210 ;
        RECT  2.075 -0.210 2.245 0.415 ;
        RECT  1.525 -0.210 2.075 0.210 ;
        RECT  1.355 -0.210 1.525 0.415 ;
        RECT  0.805 -0.210 1.355 0.210 ;
        RECT  0.635 -0.210 0.805 0.415 ;
        RECT  0.000 -0.210 0.635 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.965 2.310 11.480 2.730 ;
        RECT  2.795 1.585 2.965 2.730 ;
        RECT  2.245 2.310 2.795 2.730 ;
        RECT  2.075 1.585 2.245 2.730 ;
        RECT  1.525 2.310 2.075 2.730 ;
        RECT  1.355 1.585 1.525 2.730 ;
        RECT  0.805 2.310 1.355 2.730 ;
        RECT  0.635 1.325 0.805 2.730 ;
        RECT  0.000 2.310 0.635 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.480 2.520 ;
        LAYER M1 ;
        RECT  10.355 1.630 10.525 2.140 ;
        RECT  9.805 2.000 10.355 2.140 ;
        RECT  9.635 1.630 9.805 2.140 ;
        RECT  9.085 2.000 9.635 2.140 ;
        RECT  8.915 1.630 9.085 2.140 ;
        RECT  8.365 2.000 8.915 2.140 ;
        RECT  8.195 1.185 8.365 2.140 ;
        RECT  7.645 1.185 8.195 1.325 ;
        RECT  7.835 1.450 8.005 2.140 ;
        RECT  7.285 2.000 7.835 2.140 ;
        RECT  7.475 1.185 7.645 1.875 ;
        RECT  6.925 1.185 7.475 1.325 ;
        RECT  7.115 1.450 7.285 2.140 ;
        RECT  6.565 2.000 7.115 2.140 ;
        RECT  6.755 1.185 6.925 1.875 ;
        RECT  6.205 1.185 6.755 1.325 ;
        RECT  6.395 1.450 6.565 2.140 ;
        RECT  5.845 2.000 6.395 2.140 ;
        RECT  6.035 1.185 6.205 1.875 ;
        RECT  5.675 1.170 5.845 2.140 ;
        RECT  5.125 1.170 5.675 1.310 ;
        RECT  5.315 1.435 5.485 2.130 ;
        RECT  4.765 1.990 5.315 2.130 ;
        RECT  4.955 1.170 5.125 1.860 ;
        RECT  4.405 1.170 4.955 1.310 ;
        RECT  4.595 1.435 4.765 2.130 ;
        RECT  4.045 1.990 4.595 2.130 ;
        RECT  4.235 1.170 4.405 1.860 ;
        RECT  3.685 1.170 4.235 1.310 ;
        RECT  3.875 1.435 4.045 2.130 ;
        RECT  3.325 1.990 3.875 2.130 ;
        RECT  3.515 1.170 3.685 1.860 ;
        RECT  3.155 1.170 3.325 2.130 ;
        RECT  2.605 1.170 3.155 1.310 ;
        RECT  2.435 1.170 2.605 1.995 ;
        RECT  1.885 1.170 2.435 1.310 ;
        RECT  1.715 1.170 1.885 1.995 ;
        RECT  1.165 1.170 1.715 1.310 ;
        RECT  0.995 1.170 1.165 1.995 ;
    END
END NOR4X8AD
MACRO NOR4XLAD
    CLASS CORE ;
    FOREIGN NOR4XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 1.425 1.525 1.750 ;
        RECT  1.170 0.610 1.290 1.750 ;
        RECT  1.115 0.610 1.170 0.995 ;
        RECT  0.565 0.875 1.115 0.995 ;
        RECT  0.395 0.610 0.565 0.995 ;
        END
        AntennaDiffArea 0.205 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.590 0.230 1.285 ;
        END
        AntennaGateArea 0.064 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.115 0.760 1.375 ;
        END
        AntennaGateArea 0.064 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.115 1.050 1.650 ;
        END
        AntennaGateArea 0.064 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.465 0.605 1.610 1.285 ;
        END
        AntennaGateArea 0.064 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.515 -0.210 1.680 0.210 ;
        RECT  1.345 -0.210 1.515 0.350 ;
        RECT  0.970 -0.210 1.345 0.210 ;
        RECT  0.710 -0.210 0.970 0.755 ;
        RECT  0.335 -0.210 0.710 0.210 ;
        RECT  0.165 -0.210 0.335 0.350 ;
        RECT  0.000 -0.210 0.165 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.325 2.310 1.680 2.730 ;
        RECT  0.155 1.580 0.325 2.730 ;
        RECT  0.000 2.310 0.155 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
	 END
END NOR4XLAD
MACRO OA21X1AD
    CLASS CORE ;
    FOREIGN OA21X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.595 0.385 1.610 1.700 ;
        RECT  1.470 0.385 1.595 1.985 ;
        RECT  1.425 0.385 1.470 0.555 ;
        RECT  1.425 1.555 1.470 1.985 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 1.025 1.065 1.385 ;
        END
        AntennaGateArea 0.0414 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.205 1.045 0.375 1.375 ;
        RECT  0.070 1.145 0.205 1.375 ;
        END
        AntennaGateArea 0.041 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.495 1.025 0.770 1.375 ;
        END
        AntennaGateArea 0.041 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.235 -0.210 1.680 0.210 ;
        RECT  1.065 -0.210 1.235 0.525 ;
        RECT  0.545 -0.210 1.065 0.210 ;
        RECT  0.375 -0.210 0.545 0.905 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.215 2.310 1.680 2.730 ;
        RECT  1.045 1.935 1.215 2.730 ;
        RECT  0.255 2.310 1.045 2.730 ;
        RECT  0.085 1.495 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.185 0.735 1.305 1.625 ;
        RECT  1.045 0.735 1.185 0.905 ;
        RECT  0.915 1.505 1.185 1.625 ;
        RECT  0.850 1.505 0.915 1.675 ;
        RECT  0.730 1.505 0.850 2.185 ;
        RECT  0.680 2.015 0.730 2.185 ;
    END
END OA21X1AD
MACRO OA21X2AD
    CLASS CORE ;
    FOREIGN OA21X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.945 0.400 2.115 1.675 ;
        RECT  1.935 0.400 1.945 0.830 ;
        RECT  1.890 1.425 1.945 1.675 ;
        RECT  1.720 1.425 1.890 2.165 ;
        RECT  1.695 1.735 1.720 2.165 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.010 1.350 1.375 ;
        END
        AntennaGateArea 0.0754 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.010 0.490 1.375 ;
        END
        AntennaGateArea 0.0754 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 1.055 1.050 1.375 ;
        END
        AntennaGateArea 0.075 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.745 -0.210 2.240 0.210 ;
        RECT  1.575 -0.210 1.745 0.590 ;
        RECT  0.665 -0.210 1.575 0.210 ;
        RECT  0.495 -0.210 0.665 0.575 ;
        RECT  0.000 -0.210 0.495 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.505 2.310 2.240 2.730 ;
        RECT  1.335 1.785 1.505 2.730 ;
        RECT  0.385 2.310 1.335 2.730 ;
        RECT  0.215 1.495 0.385 2.730 ;
        RECT  0.000 2.310 0.215 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.600 1.065 1.745 1.235 ;
        RECT  1.480 0.770 1.600 1.615 ;
        RECT  1.405 0.770 1.480 0.890 ;
        RECT  1.045 1.495 1.480 1.615 ;
        RECT  1.235 0.680 1.405 0.890 ;
        RECT  0.115 0.695 1.045 0.865 ;
        RECT  0.875 1.495 1.045 1.665 ;
    END
END OA21X2AD
MACRO OA21X4AD
    CLASS CORE ;
    FOREIGN OA21X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.045 1.005 2.170 1.515 ;
        RECT  1.875 0.385 2.045 1.515 ;
        RECT  1.725 1.345 1.875 1.515 ;
        RECT  1.555 1.345 1.725 1.960 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.065 1.125 1.375 ;
        END
        AntennaGateArea 0.1455 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.205 1.055 0.435 1.375 ;
        RECT  0.070 1.140 0.205 1.375 ;
        END
        AntennaGateArea 0.144 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 1.045 0.790 1.375 ;
        END
        AntennaGateArea 0.144 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.405 -0.210 2.520 0.210 ;
        RECT  2.235 -0.210 2.405 0.815 ;
        RECT  1.685 -0.210 2.235 0.210 ;
        RECT  1.515 -0.210 1.685 0.815 ;
        RECT  0.640 -0.210 1.515 0.210 ;
        RECT  0.420 -0.210 0.640 0.595 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.085 2.310 2.520 2.730 ;
        RECT  1.915 1.635 2.085 2.730 ;
        RECT  1.365 2.310 1.915 2.730 ;
        RECT  1.195 1.735 1.365 2.730 ;
        RECT  0.315 2.310 1.195 2.730 ;
        RECT  0.145 1.495 0.315 2.730 ;
        RECT  0.000 2.310 0.145 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.385 1.055 1.745 1.225 ;
        RECT  1.335 0.795 1.385 1.615 ;
        RECT  1.245 0.415 1.335 1.615 ;
        RECT  1.165 0.415 1.245 0.915 ;
        RECT  0.975 1.495 1.245 1.615 ;
        RECT  0.805 0.390 0.975 0.920 ;
        RECT  0.805 1.495 0.975 1.925 ;
        RECT  0.255 0.760 0.805 0.920 ;
        RECT  0.085 0.390 0.255 0.920 ;
    END
END OA21X4AD
MACRO OA21XLAD
    CLASS CORE ;
    FOREIGN OA21XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.385 1.610 1.865 ;
        RECT  1.425 0.385 1.470 0.555 ;
        RECT  1.425 1.695 1.470 1.865 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 1.025 1.065 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.205 1.045 0.375 1.375 ;
        RECT  0.070 1.145 0.205 1.375 ;
        END
        AntennaGateArea 0.04 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.495 1.025 0.770 1.375 ;
        END
        AntennaGateArea 0.04 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.235 -0.210 1.680 0.210 ;
        RECT  1.065 -0.210 1.235 0.555 ;
        RECT  0.545 -0.210 1.065 0.210 ;
        RECT  0.375 -0.210 0.545 0.905 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.215 2.310 1.680 2.730 ;
        RECT  1.045 1.925 1.215 2.730 ;
        RECT  0.255 2.310 1.045 2.730 ;
        RECT  0.085 1.495 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.185 0.735 1.305 1.615 ;
        RECT  1.045 0.735 1.185 0.905 ;
        RECT  0.915 1.495 1.185 1.615 ;
        RECT  0.850 1.495 0.915 1.665 ;
        RECT  0.730 1.495 0.850 2.185 ;
        RECT  0.680 2.015 0.730 2.185 ;
    END
END OA21XLAD
MACRO OA22X1AD
    CLASS CORE ;
    FOREIGN OA22X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.155 0.430 2.170 1.555 ;
        RECT  2.010 0.385 2.155 1.805 ;
        RECT  1.985 0.385 2.010 0.555 ;
        RECT  1.985 1.375 2.010 1.805 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 0.820 1.640 1.250 ;
        RECT  1.470 0.820 1.610 1.375 ;
        END
        AntennaGateArea 0.0464 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.070 1.330 1.375 ;
        RECT  1.030 1.050 1.150 1.375 ;
        RECT  1.000 1.070 1.030 1.375 ;
        END
        AntennaGateArea 0.046 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.225 1.080 0.270 1.300 ;
        RECT  0.210 1.060 0.225 1.320 ;
        RECT  0.105 1.060 0.210 1.655 ;
        RECT  0.070 1.080 0.105 1.655 ;
        END
        AntennaGateArea 0.0464 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.025 0.870 1.375 ;
        END
        AntennaGateArea 0.046 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.795 -0.210 2.240 0.210 ;
        RECT  1.625 -0.210 1.795 0.555 ;
        RECT  1.055 -0.210 1.625 0.210 ;
        RECT  0.885 -0.210 1.055 0.375 ;
        RECT  0.000 -0.210 0.885 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.795 2.310 2.240 2.730 ;
        RECT  1.625 1.525 1.795 2.730 ;
        RECT  0.265 2.310 1.625 2.730 ;
        RECT  0.095 1.775 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.355 2.005 1.480 2.175 ;
        RECT  1.345 0.385 1.435 0.555 ;
        RECT  1.235 1.500 1.355 2.175 ;
        RECT  1.225 0.385 1.345 0.905 ;
        RECT  0.510 1.500 1.235 1.620 ;
        RECT  0.975 0.785 1.225 0.905 ;
        RECT  0.905 0.735 0.975 0.905 ;
        RECT  0.785 0.495 0.905 0.905 ;
        RECT  0.255 0.495 0.785 0.615 ;
        RECT  0.510 0.735 0.615 0.905 ;
        RECT  0.390 0.735 0.510 1.620 ;
        RECT  0.135 0.495 0.255 0.905 ;
        RECT  0.085 0.735 0.135 0.905 ;
    END
END OA22X1AD
MACRO OA22X2AD
    CLASS CORE ;
    FOREIGN OA22X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.435 0.680 2.450 2.035 ;
        RECT  2.290 0.395 2.435 2.035 ;
        RECT  2.265 0.395 2.290 0.825 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.115 1.845 1.375 ;
        END
        AntennaGateArea 0.0843 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.095 1.350 1.375 ;
        END
        AntennaGateArea 0.084 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.225 1.140 0.270 1.360 ;
        RECT  0.210 1.120 0.225 1.380 ;
        RECT  0.105 1.120 0.210 1.655 ;
        RECT  0.070 1.140 0.105 1.655 ;
        END
        AntennaGateArea 0.0853 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.095 0.910 1.375 ;
        END
        AntennaGateArea 0.084 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.055 -0.210 2.520 0.210 ;
        RECT  2.055 0.395 2.065 0.825 ;
        RECT  1.895 -0.210 2.055 0.825 ;
        RECT  1.885 -0.210 1.895 0.560 ;
        RECT  1.325 -0.210 1.885 0.210 ;
        RECT  1.155 -0.210 1.325 0.735 ;
        RECT  0.000 -0.210 1.155 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.945 2.310 2.520 2.730 ;
        RECT  1.775 1.735 1.945 2.730 ;
        RECT  0.295 2.310 1.775 2.730 ;
        RECT  0.125 1.775 0.295 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.115 1.065 2.165 1.235 ;
        RECT  1.995 1.065 2.115 1.615 ;
        RECT  1.235 1.495 1.995 1.615 ;
        RECT  1.635 0.675 1.685 0.845 ;
        RECT  1.515 0.675 1.635 0.975 ;
        RECT  0.950 0.855 1.515 0.975 ;
        RECT  0.805 1.495 1.235 1.720 ;
        RECT  0.830 0.445 0.950 0.975 ;
        RECT  0.255 0.445 0.830 0.565 ;
        RECT  0.510 1.495 0.805 1.615 ;
        RECT  0.510 0.685 0.615 0.855 ;
        RECT  0.390 0.685 0.510 1.615 ;
        RECT  0.135 0.445 0.255 0.815 ;
        RECT  0.085 0.645 0.135 0.815 ;
    END
END OA22X2AD
MACRO OA22X4AD
    CLASS CORE ;
    FOREIGN OA22X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.705 1.285 2.730 1.990 ;
        RECT  2.575 0.360 2.705 1.990 ;
        RECT  2.465 0.360 2.575 0.790 ;
        RECT  2.465 1.560 2.575 1.990 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.050 2.010 1.375 ;
        RECT  1.730 1.110 1.750 1.230 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.020 1.610 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.065 0.440 1.375 ;
        RECT  0.070 1.145 0.210 1.655 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 1.020 1.150 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.995 -0.210 3.080 0.210 ;
        RECT  2.825 -0.210 2.995 0.815 ;
        RECT  2.235 -0.210 2.825 0.210 ;
        RECT  2.065 -0.210 2.235 0.795 ;
        RECT  1.480 -0.210 2.065 0.210 ;
        RECT  1.220 -0.210 1.480 0.650 ;
        RECT  0.000 -0.210 1.220 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.980 2.310 3.080 2.730 ;
        RECT  2.850 1.495 2.980 2.730 ;
        RECT  2.160 2.310 2.850 2.730 ;
        RECT  1.990 1.845 2.160 2.730 ;
        RECT  0.355 2.310 1.990 2.730 ;
        RECT  0.185 1.845 0.355 2.730 ;
        RECT  0.000 2.310 0.185 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  2.250 1.065 2.455 1.235 ;
        RECT  2.130 1.065 2.250 1.705 ;
        RECT  1.335 1.495 2.130 1.705 ;
        RECT  1.645 0.360 1.815 0.900 ;
        RECT  1.015 0.780 1.645 0.900 ;
        RECT  0.905 1.495 1.335 1.970 ;
        RECT  0.845 0.390 1.015 0.900 ;
        RECT  0.680 1.495 0.905 1.705 ;
        RECT  0.295 0.390 0.845 0.510 ;
        RECT  0.560 0.630 0.680 1.705 ;
        RECT  0.485 0.630 0.560 0.800 ;
        RECT  0.125 0.390 0.295 0.820 ;
    END
END OA22X4AD
MACRO OA22XLAD
    CLASS CORE ;
    FOREIGN OA22XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.385 2.170 1.675 ;
        RECT  1.985 0.385 2.030 0.555 ;
        RECT  1.985 1.505 2.030 1.675 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 0.820 1.640 1.250 ;
        RECT  1.470 0.820 1.610 1.375 ;
        END
        AntennaGateArea 0.04 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.070 1.330 1.375 ;
        RECT  1.030 1.050 1.150 1.375 ;
        RECT  1.000 1.070 1.030 1.375 ;
        END
        AntennaGateArea 0.04 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.225 1.080 0.270 1.300 ;
        RECT  0.210 1.060 0.225 1.320 ;
        RECT  0.105 1.060 0.210 1.655 ;
        RECT  0.070 1.080 0.105 1.655 ;
        END
        AntennaGateArea 0.0404 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.025 0.870 1.375 ;
        END
        AntennaGateArea 0.04 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.795 -0.210 2.240 0.210 ;
        RECT  1.625 -0.210 1.795 0.555 ;
        RECT  1.055 -0.210 1.625 0.210 ;
        RECT  0.885 -0.210 1.055 0.375 ;
        RECT  0.000 -0.210 0.885 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.795 2.310 2.240 2.730 ;
        RECT  1.625 1.505 1.795 2.730 ;
        RECT  0.265 2.310 1.625 2.730 ;
        RECT  0.095 1.775 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.355 2.005 1.480 2.175 ;
        RECT  1.345 0.385 1.435 0.555 ;
        RECT  1.235 1.500 1.355 2.175 ;
        RECT  1.225 0.385 1.345 0.905 ;
        RECT  0.510 1.500 1.235 1.620 ;
        RECT  0.975 0.785 1.225 0.905 ;
        RECT  0.905 0.735 0.975 0.905 ;
        RECT  0.785 0.495 0.905 0.905 ;
        RECT  0.255 0.495 0.785 0.615 ;
        RECT  0.510 0.735 0.615 0.905 ;
        RECT  0.390 0.735 0.510 1.620 ;
        RECT  0.135 0.495 0.255 0.905 ;
        RECT  0.085 0.735 0.135 0.905 ;
    END
END OA22XLAD
MACRO OAI211X1AD
    CLASS CORE ;
    FOREIGN OAI211X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.570 0.645 1.610 1.655 ;
        RECT  1.450 0.645 1.570 1.935 ;
        RECT  0.895 1.495 1.450 1.655 ;
        RECT  0.725 1.495 0.895 1.925 ;
        END
        AntennaDiffArea 0.36 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.025 1.070 1.375 ;
        END
        AntennaGateArea 0.0884 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 0.335 1.475 0.505 ;
        RECT  1.190 0.335 1.330 1.375 ;
        END
        AntennaGateArea 0.0884 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.025 0.230 1.655 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 1.025 0.720 1.285 ;
        RECT  0.600 1.025 0.685 1.290 ;
        RECT  0.490 1.070 0.600 1.290 ;
        RECT  0.350 1.070 0.490 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.680 -0.210 1.680 0.210 ;
        RECT  0.420 -0.210 0.680 0.360 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.310 1.680 2.730 ;
        RECT  1.240 2.230 1.260 2.730 ;
        RECT  1.020 2.185 1.240 2.730 ;
        RECT  1.000 2.230 1.020 2.730 ;
        RECT  0.285 2.310 1.000 2.730 ;
        RECT  0.115 1.780 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  0.815 0.710 0.985 0.880 ;
        RECT  0.255 0.760 0.815 0.880 ;
        RECT  0.085 0.710 0.255 0.880 ;
    END
END OAI211X1AD
MACRO OAI211X2AD
    CLASS CORE ;
    FOREIGN OAI211X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.740 1.890 1.720 ;
        RECT  1.645 0.740 1.750 0.880 ;
        RECT  1.685 1.550 1.750 1.720 ;
        RECT  1.515 1.550 1.685 1.980 ;
        RECT  1.475 0.405 1.645 0.880 ;
        RECT  0.925 1.550 1.515 1.720 ;
        RECT  0.755 1.550 0.925 1.980 ;
        END
        AntennaDiffArea 0.615 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 1.055 1.170 1.430 ;
        END
        AntennaGateArea 0.162 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.000 1.630 1.430 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 1.065 0.385 1.235 ;
        RECT  0.070 1.065 0.230 1.655 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.525 1.055 0.770 1.430 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.625 -0.210 1.960 0.210 ;
        RECT  0.455 -0.210 0.625 0.675 ;
        RECT  0.000 -0.210 0.455 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.305 2.310 1.960 2.730 ;
        RECT  1.135 1.845 1.305 2.730 ;
        RECT  0.265 2.310 1.135 2.730 ;
        RECT  0.095 1.845 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  0.815 0.405 0.985 0.915 ;
        RECT  0.265 0.795 0.815 0.915 ;
        RECT  0.095 0.405 0.265 0.915 ;
    END
END OAI211X2AD
MACRO OAI211X4AD
    CLASS CORE ;
    FOREIGN OAI211X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.135 0.785 3.155 1.660 ;
        RECT  3.025 0.785 3.135 1.960 ;
        RECT  2.735 0.785 3.025 0.915 ;
        RECT  2.965 1.530 3.025 1.960 ;
        RECT  2.415 1.530 2.965 1.660 ;
        RECT  2.615 0.670 2.735 0.915 ;
        RECT  2.200 0.670 2.615 0.790 ;
        RECT  2.245 1.530 2.415 1.980 ;
        RECT  1.675 1.530 2.245 1.660 ;
        RECT  1.460 1.530 1.675 2.085 ;
        RECT  0.335 1.530 1.460 1.660 ;
        RECT  0.325 1.530 0.335 1.760 ;
        RECT  0.155 1.530 0.325 1.960 ;
        END
        AntennaDiffArea 1.092 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.780 1.035 2.900 1.410 ;
        RECT  1.935 1.290 2.780 1.410 ;
        RECT  1.815 0.910 1.935 1.410 ;
        RECT  1.740 0.910 1.815 1.260 ;
        RECT  1.705 0.910 1.740 1.240 ;
        END
        AntennaGateArea 0.324 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.110 0.910 2.495 1.170 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.120 1.190 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 0.880 1.500 1.280 ;
        RECT  0.535 0.880 1.380 1.000 ;
        RECT  0.450 0.880 0.535 1.235 ;
        RECT  0.330 0.880 0.450 1.255 ;
        RECT  0.305 0.880 0.330 1.235 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.395 -0.210 3.360 0.210 ;
        RECT  1.225 -0.210 1.395 0.485 ;
        RECT  0.625 -0.210 1.225 0.210 ;
        RECT  0.455 -0.210 0.625 0.485 ;
        RECT  0.000 -0.210 0.455 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.775 2.310 3.360 2.730 ;
        RECT  2.605 1.845 2.775 2.730 ;
        RECT  2.005 2.310 2.605 2.730 ;
        RECT  1.835 1.845 2.005 2.730 ;
        RECT  0.985 2.310 1.835 2.730 ;
        RECT  0.815 1.845 0.985 2.730 ;
        RECT  0.000 2.310 0.815 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  1.755 0.430 3.120 0.550 ;
        RECT  1.585 0.330 1.755 0.760 ;
        RECT  0.985 0.640 1.585 0.760 ;
        RECT  0.815 0.330 0.985 0.760 ;
        RECT  0.265 0.640 0.815 0.760 ;
        RECT  0.095 0.330 0.265 0.760 ;
    END
END OAI211X4AD
MACRO OAI211XLAD
    CLASS CORE ;
    FOREIGN OAI211XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 0.690 1.610 1.655 ;
        RECT  0.895 1.495 1.450 1.655 ;
        RECT  0.725 1.495 0.895 1.665 ;
        END
        AntennaDiffArea 0.242 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.025 1.070 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 0.400 1.475 0.570 ;
        RECT  1.190 0.400 1.330 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.025 0.230 1.460 ;
        END
        AntennaGateArea 0.06 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 1.025 0.720 1.285 ;
        RECT  0.600 1.025 0.685 1.290 ;
        RECT  0.490 1.070 0.600 1.290 ;
        RECT  0.350 1.070 0.490 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.680 -0.210 1.680 0.210 ;
        RECT  0.420 -0.210 0.680 0.540 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.215 2.310 1.680 2.730 ;
        RECT  1.045 1.995 1.215 2.730 ;
        RECT  0.285 2.310 1.045 2.730 ;
        RECT  0.115 1.580 0.285 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  0.815 0.735 0.985 0.905 ;
        RECT  0.255 0.785 0.815 0.905 ;
        RECT  0.085 0.735 0.255 0.905 ;
    END
END OAI211XLAD
MACRO OAI21BX1AD
    CLASS CORE ;
    FOREIGN OAI21BX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.385 1.275 0.555 ;
        RECT  0.925 0.385 1.050 1.665 ;
        RECT  0.910 0.385 0.925 1.955 ;
        RECT  0.755 1.525 0.910 1.955 ;
        END
        AntennaDiffArea 0.257 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.585 1.890 1.200 ;
        RECT  1.420 1.080 1.750 1.200 ;
        END
        AntennaGateArea 0.0414 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.270 1.030 0.390 1.375 ;
        RECT  0.070 1.145 0.270 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 0.955 0.770 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.835 -0.210 1.960 0.210 ;
        RECT  1.575 -0.210 1.835 0.450 ;
        RECT  0.545 -0.210 1.575 0.210 ;
        RECT  0.375 -0.210 0.545 0.815 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.430 2.310 1.960 2.730 ;
        RECT  1.170 1.560 1.430 2.730 ;
        RECT  0.265 2.310 1.170 2.730 ;
        RECT  0.095 1.525 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.605 1.320 1.775 1.555 ;
        RECT  1.290 1.320 1.605 1.440 ;
        RECT  1.390 0.690 1.510 0.950 ;
        RECT  1.290 0.830 1.390 0.950 ;
        RECT  1.170 0.830 1.290 1.440 ;
    END
END OAI21BX1AD
MACRO OAI21BX2AD
    CLASS CORE ;
    FOREIGN OAI21BX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.310 0.385 1.425 0.815 ;
        RECT  1.190 0.385 1.310 1.000 ;
        RECT  1.125 0.880 1.190 1.000 ;
        RECT  1.005 0.880 1.125 1.975 ;
        RECT  0.885 1.545 1.005 1.975 ;
        END
        AntennaDiffArea 0.425 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.865 2.170 1.390 ;
        RECT  1.845 1.025 2.030 1.195 ;
        END
        AntennaGateArea 0.065 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.365 1.040 0.510 1.375 ;
        RECT  0.070 1.145 0.365 1.375 ;
        END
        AntennaGateArea 0.1629 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.040 0.865 1.415 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.135 -0.210 2.240 0.210 ;
        RECT  1.965 -0.210 2.135 0.745 ;
        RECT  0.665 -0.210 1.965 0.210 ;
        RECT  0.495 -0.210 0.665 0.485 ;
        RECT  0.000 -0.210 0.495 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.435 2.310 2.240 2.730 ;
        RECT  1.265 1.560 1.435 2.730 ;
        RECT  0.380 2.310 1.265 2.730 ;
        RECT  0.210 1.600 0.380 2.730 ;
        RECT  0.000 2.310 0.210 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.770 1.510 1.940 1.680 ;
        RECT  1.725 0.610 1.775 0.780 ;
        RECT  1.725 1.510 1.770 1.630 ;
        RECT  1.605 0.610 1.725 1.630 ;
        RECT  1.245 1.120 1.605 1.240 ;
        RECT  0.885 0.330 1.055 0.760 ;
        RECT  0.290 0.640 0.885 0.760 ;
        RECT  0.120 0.330 0.290 0.760 ;
    END
END OAI21BX2AD
MACRO OAI21BX4AD
    CLASS CORE ;
    FOREIGN OAI21BX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.900 0.730 2.070 1.990 ;
        RECT  1.750 1.005 1.900 1.580 ;
        RECT  0.990 1.450 1.750 1.580 ;
        RECT  0.820 1.450 0.990 2.010 ;
        END
        AntennaDiffArea 0.664 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.100 1.145 3.290 1.375 ;
        RECT  2.980 1.020 3.100 1.540 ;
        END
        AntennaGateArea 0.1295 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.355 0.900 1.475 1.260 ;
        RECT  0.650 0.900 1.355 1.020 ;
        RECT  0.530 0.900 0.650 1.140 ;
        RECT  0.490 1.020 0.530 1.140 ;
        RECT  0.335 1.020 0.490 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.140 1.160 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.180 -0.210 3.360 0.210 ;
        RECT  3.010 -0.210 3.180 0.745 ;
        RECT  1.350 -0.210 3.010 0.210 ;
        RECT  1.180 -0.210 1.350 0.470 ;
        RECT  0.630 -0.210 1.180 0.210 ;
        RECT  0.460 -0.210 0.630 0.470 ;
        RECT  0.000 -0.210 0.460 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.430 2.310 3.360 2.730 ;
        RECT  2.260 1.665 2.430 2.730 ;
        RECT  1.655 2.310 2.260 2.730 ;
        RECT  1.485 1.735 1.655 2.730 ;
        RECT  0.330 2.310 1.485 2.730 ;
        RECT  0.160 1.735 0.330 2.730 ;
        RECT  0.000 2.310 0.160 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.790 1.385 2.840 1.890 ;
        RECT  2.670 0.475 2.790 1.890 ;
        RECT  2.620 0.475 2.670 1.555 ;
        RECT  2.190 1.065 2.620 1.235 ;
        RECT  2.260 0.350 2.430 0.780 ;
        RECT  1.710 0.440 2.260 0.610 ;
        RECT  1.540 0.350 1.710 0.780 ;
        RECT  0.990 0.660 1.540 0.780 ;
        RECT  0.820 0.350 0.990 0.780 ;
        RECT  0.270 0.660 0.820 0.780 ;
        RECT  0.100 0.350 0.270 0.780 ;
    END
END OAI21BX4AD
MACRO OAI21BXLAD
    CLASS CORE ;
    FOREIGN OAI21BXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.385 1.275 0.555 ;
        RECT  0.925 0.385 1.050 1.665 ;
        RECT  0.910 0.385 0.925 1.695 ;
        RECT  0.755 1.525 0.910 1.695 ;
        END
        AntennaDiffArea 0.198 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.585 1.890 1.200 ;
        RECT  1.420 1.080 1.750 1.200 ;
        END
        AntennaGateArea 0.0403 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.270 1.030 0.390 1.375 ;
        RECT  0.070 1.145 0.270 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 1.025 0.770 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.790 -0.210 1.960 0.210 ;
        RECT  1.620 -0.210 1.790 0.465 ;
        RECT  0.545 -0.210 1.620 0.210 ;
        RECT  0.375 -0.210 0.545 0.905 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.430 2.310 1.960 2.730 ;
        RECT  1.170 1.560 1.430 2.730 ;
        RECT  0.265 2.310 1.170 2.730 ;
        RECT  0.095 1.525 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.605 1.320 1.775 1.555 ;
        RECT  1.290 1.320 1.605 1.440 ;
        RECT  1.390 0.690 1.510 0.950 ;
        RECT  1.290 0.830 1.390 0.950 ;
        RECT  1.170 0.830 1.290 1.440 ;
    END
END OAI21BXLAD
MACRO OAI21X1AD
    CLASS CORE ;
    FOREIGN OAI21X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.695 1.330 1.665 ;
        RECT  1.135 0.695 1.190 0.865 ;
        RECT  0.980 1.545 1.190 1.665 ;
        RECT  0.720 1.545 0.980 1.925 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 1.030 1.070 1.425 ;
        RECT  0.925 1.010 1.045 1.425 ;
        RECT  0.900 1.030 0.925 1.425 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.280 1.020 0.400 1.375 ;
        RECT  0.070 1.145 0.280 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.020 0.770 1.425 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.565 -0.210 1.400 0.210 ;
        RECT  0.395 -0.210 0.565 0.385 ;
        RECT  0.000 -0.210 0.395 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.295 2.310 1.400 2.730 ;
        RECT  1.125 1.785 1.295 2.730 ;
        RECT  0.275 2.310 1.125 2.730 ;
        RECT  0.105 1.495 0.275 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.085 0.695 0.945 0.865 ;
    END
END OAI21X1AD
MACRO OAI21X2AD
    CLASS CORE ;
    FOREIGN OAI21X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.520 0.685 1.610 1.625 ;
        RECT  1.470 0.400 1.520 1.625 ;
        RECT  1.350 0.400 1.470 0.830 ;
        RECT  1.040 1.495 1.470 1.625 ;
        RECT  0.870 1.495 1.040 2.035 ;
        END
        AntennaDiffArea 0.457 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.040 1.260 1.375 ;
        END
        AntennaGateArea 0.1629 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 1.040 0.440 1.375 ;
        RECT  0.210 1.145 0.320 1.375 ;
        RECT  0.070 1.145 0.210 1.655 ;
        END
        AntennaGateArea 0.1629 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 1.035 0.790 1.375 ;
        END
        AntennaGateArea 0.1629 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.740 -0.210 1.680 0.210 ;
        RECT  0.570 -0.210 0.740 0.675 ;
        RECT  0.000 -0.210 0.570 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.430 2.310 1.680 2.730 ;
        RECT  1.260 1.775 1.430 2.730 ;
        RECT  0.350 2.310 1.260 2.730 ;
        RECT  0.180 1.775 0.350 2.730 ;
        RECT  0.000 2.310 0.180 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  0.980 0.400 1.150 0.915 ;
        RECT  0.350 0.795 0.980 0.915 ;
        RECT  0.180 0.400 0.350 0.915 ;
    END
END OAI21X2AD
MACRO OAI21X3AD
    CLASS CORE ;
    FOREIGN OAI21X3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.055 0.690 2.170 1.795 ;
        RECT  2.030 0.690 2.055 1.925 ;
        RECT  1.885 0.690 2.030 0.860 ;
        RECT  1.885 1.495 2.030 1.925 ;
        RECT  0.975 1.495 1.885 1.665 ;
        RECT  0.805 1.495 0.975 1.925 ;
        END
        AntennaDiffArea 0.5 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.880 1.030 1.905 1.375 ;
        RECT  1.760 1.020 1.880 1.375 ;
        RECT  1.605 1.030 1.760 1.375 ;
        END
        AntennaGateArea 0.244 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 0.900 1.460 1.280 ;
        RECT  0.460 0.900 1.340 1.020 ;
        RECT  0.340 0.900 0.460 1.375 ;
        RECT  0.320 1.020 0.340 1.375 ;
        RECT  0.070 1.145 0.320 1.375 ;
        END
        AntennaGateArea 0.244 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.110 1.140 1.140 1.260 ;
        RECT  0.630 1.140 1.110 1.375 ;
        RECT  0.620 1.140 0.630 1.260 ;
        END
        AntennaGateArea 0.2447 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.335 -0.210 2.520 0.210 ;
        RECT  1.165 -0.210 1.335 0.540 ;
        RECT  0.615 -0.210 1.165 0.210 ;
        RECT  0.445 -0.210 0.615 0.540 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 2.310 2.520 2.730 ;
        RECT  2.290 1.510 2.410 2.730 ;
        RECT  1.635 2.310 2.290 2.730 ;
        RECT  1.465 1.825 1.635 2.730 ;
        RECT  0.315 2.310 1.465 2.730 ;
        RECT  0.145 1.555 0.315 2.730 ;
        RECT  0.000 2.310 0.145 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.290 0.385 2.410 0.905 ;
        RECT  1.740 0.450 2.290 0.570 ;
        RECT  1.480 0.400 1.740 0.780 ;
        RECT  1.020 0.660 1.480 0.780 ;
        RECT  0.760 0.400 1.020 0.780 ;
        RECT  0.255 0.660 0.760 0.780 ;
        RECT  0.085 0.375 0.255 0.805 ;
    END
END OAI21X3AD
MACRO OAI21X4AD
    CLASS CORE ;
    FOREIGN OAI21X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.055 0.755 2.170 1.795 ;
        RECT  2.030 0.725 2.055 2.005 ;
        RECT  1.885 0.725 2.030 0.895 ;
        RECT  1.885 1.555 2.030 2.005 ;
        RECT  0.975 1.555 1.885 1.725 ;
        RECT  0.805 1.555 0.975 2.005 ;
        END
        AntennaDiffArea 0.664 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.655 1.015 1.905 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 0.870 1.460 1.280 ;
        RECT  0.440 0.870 1.340 0.990 ;
        RECT  0.320 0.870 0.440 1.375 ;
        RECT  0.070 1.145 0.320 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.110 1.150 1.380 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.335 -0.210 2.520 0.210 ;
        RECT  1.165 -0.210 1.335 0.510 ;
        RECT  0.615 -0.210 1.165 0.210 ;
        RECT  0.445 -0.210 0.615 0.510 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 2.310 2.520 2.730 ;
        RECT  2.290 1.575 2.410 2.730 ;
        RECT  1.635 2.310 2.290 2.730 ;
        RECT  1.465 1.845 1.635 2.730 ;
        RECT  0.315 2.310 1.465 2.730 ;
        RECT  0.145 1.560 0.315 2.730 ;
        RECT  0.000 2.310 0.145 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.290 0.380 2.410 0.900 ;
        RECT  1.740 0.380 2.290 0.550 ;
        RECT  1.480 0.340 1.740 0.750 ;
        RECT  1.020 0.630 1.480 0.750 ;
        RECT  0.760 0.370 1.020 0.750 ;
        RECT  0.255 0.630 0.760 0.750 ;
        RECT  0.085 0.330 0.255 0.760 ;
    END
END OAI21X4AD
MACRO OAI21X6AD
    CLASS CORE ;
    FOREIGN OAI21X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.535 0.700 3.570 1.725 ;
        RECT  3.520 0.700 3.535 1.980 ;
        RECT  3.400 0.370 3.520 1.980 ;
        RECT  2.570 0.700 3.400 0.820 ;
        RECT  3.365 1.545 3.400 1.980 ;
        RECT  2.785 1.545 3.365 1.725 ;
        RECT  2.615 1.545 2.785 1.980 ;
        RECT  1.705 1.545 2.615 1.725 ;
        RECT  1.535 1.545 1.705 1.980 ;
        RECT  0.265 1.545 1.535 1.725 ;
        RECT  0.095 1.545 0.265 1.980 ;
        END
        AntennaDiffArea 1.258 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.730 1.110 3.275 1.230 ;
        RECT  2.495 1.110 2.730 1.375 ;
        END
        AntennaGateArea 0.486 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.070 0.900 2.190 1.280 ;
        RECT  1.210 0.900 2.070 1.020 ;
        RECT  0.690 0.900 1.210 1.140 ;
        END
        AntennaGateArea 0.486 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.140 1.890 1.280 ;
        RECT  1.370 1.140 1.610 1.400 ;
        RECT  0.400 1.260 1.370 1.400 ;
        RECT  0.260 1.020 0.400 1.400 ;
        END
        AntennaGateArea 0.4869 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.065 -0.210 3.640 0.210 ;
        RECT  1.895 -0.210 2.065 0.500 ;
        RECT  1.345 -0.210 1.895 0.210 ;
        RECT  1.175 -0.210 1.345 0.500 ;
        RECT  0.625 -0.210 1.175 0.210 ;
        RECT  0.455 -0.210 0.625 0.500 ;
        RECT  0.000 -0.210 0.455 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.145 2.310 3.640 2.730 ;
        RECT  2.975 1.845 3.145 2.730 ;
        RECT  2.425 2.310 2.975 2.730 ;
        RECT  2.255 1.845 2.425 2.730 ;
        RECT  0.930 2.310 2.255 2.730 ;
        RECT  0.760 1.845 0.930 2.730 ;
        RECT  0.000 2.310 0.760 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  2.425 0.390 3.145 0.560 ;
        RECT  2.255 0.350 2.425 0.780 ;
        RECT  1.705 0.660 2.255 0.780 ;
        RECT  1.535 0.350 1.705 0.780 ;
        RECT  0.985 0.660 1.535 0.780 ;
        RECT  0.815 0.350 0.985 0.780 ;
        RECT  0.265 0.660 0.815 0.780 ;
        RECT  0.095 0.350 0.265 0.780 ;
    END
END OAI21X6AD
MACRO OAI21X8AD
    CLASS CORE ;
    FOREIGN OAI21X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.245 0.720 4.270 1.860 ;
        RECT  4.075 0.720 4.245 2.075 ;
        RECT  3.850 0.720 4.075 1.860 ;
        RECT  3.355 0.720 3.850 0.970 ;
        RECT  3.525 1.610 3.850 1.860 ;
        RECT  3.355 1.610 3.525 2.040 ;
        RECT  2.445 1.610 3.355 1.860 ;
        RECT  2.275 1.610 2.445 2.040 ;
        RECT  1.005 1.610 2.275 1.860 ;
        RECT  0.835 1.610 1.005 2.040 ;
        END
        AntennaDiffArea 1.346 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.090 3.710 1.375 ;
        END
        AntennaGateArea 0.648 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.810 0.860 2.930 1.280 ;
        RECT  1.850 0.860 2.810 0.980 ;
        RECT  1.330 0.860 1.850 1.170 ;
        RECT  0.500 0.860 1.330 0.980 ;
        RECT  0.380 0.860 0.500 1.240 ;
        END
        AntennaGateArea 0.648 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 1.100 2.610 1.240 ;
        RECT  2.230 1.100 2.450 1.375 ;
        RECT  2.090 1.100 2.230 1.430 ;
        RECT  1.170 1.290 2.090 1.430 ;
        RECT  1.030 1.100 1.170 1.430 ;
        RECT  0.650 1.100 1.030 1.220 ;
        END
        AntennaGateArea 0.648 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.805 -0.210 4.760 0.210 ;
        RECT  2.635 -0.210 2.805 0.500 ;
        RECT  2.085 -0.210 2.635 0.210 ;
        RECT  1.915 -0.210 2.085 0.500 ;
        RECT  1.365 -0.210 1.915 0.210 ;
        RECT  1.195 -0.210 1.365 0.500 ;
        RECT  0.625 -0.210 1.195 0.210 ;
        RECT  0.455 -0.210 0.625 0.500 ;
        RECT  0.000 -0.210 0.455 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.605 2.310 4.760 2.730 ;
        RECT  4.435 1.600 4.605 2.730 ;
        RECT  3.885 2.310 4.435 2.730 ;
        RECT  3.715 2.045 3.885 2.730 ;
        RECT  3.110 2.310 3.715 2.730 ;
        RECT  2.940 2.045 3.110 2.730 ;
        RECT  1.670 2.310 2.940 2.730 ;
        RECT  1.500 2.045 1.670 2.730 ;
        RECT  0.345 2.310 1.500 2.730 ;
        RECT  0.175 1.605 0.345 2.730 ;
        RECT  0.000 2.310 0.175 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.760 2.520 ;
        LAYER M1 ;
        RECT  4.460 0.380 4.580 0.900 ;
        RECT  3.210 0.380 4.460 0.550 ;
        RECT  2.950 0.360 3.210 0.740 ;
        RECT  2.490 0.620 2.950 0.740 ;
        RECT  2.230 0.360 2.490 0.740 ;
        RECT  1.770 0.620 2.230 0.740 ;
        RECT  1.510 0.360 1.770 0.740 ;
        RECT  1.040 0.620 1.510 0.740 ;
        RECT  0.780 0.360 1.040 0.740 ;
        RECT  0.265 0.620 0.780 0.740 ;
        RECT  0.095 0.330 0.265 0.760 ;
    END
END OAI21X8AD
MACRO OAI21XLAD
    CLASS CORE ;
    FOREIGN OAI21XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.305 0.735 1.330 1.665 ;
        RECT  1.190 0.730 1.305 1.665 ;
        RECT  1.135 0.730 1.190 0.900 ;
        RECT  0.720 1.545 1.190 1.665 ;
        END
        AntennaDiffArea 0.15 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.900 1.020 1.070 1.425 ;
        END
        AntennaGateArea 0.0604 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.280 1.020 0.400 1.375 ;
        RECT  0.070 1.145 0.280 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.020 0.770 1.425 ;
        END
        AntennaGateArea 0.06 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.565 -0.210 1.400 0.210 ;
        RECT  0.395 -0.210 0.565 0.470 ;
        RECT  0.000 -0.210 0.395 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.315 2.310 1.400 2.730 ;
        RECT  1.145 1.785 1.315 2.730 ;
        RECT  0.275 2.310 1.145 2.730 ;
        RECT  0.105 1.495 0.275 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.085 0.730 0.945 0.900 ;
    END
END OAI21XLAD
MACRO OAI221X1AD
    CLASS CORE ;
    FOREIGN OAI221X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.365 0.705 2.450 1.655 ;
        RECT  2.310 0.705 2.365 1.945 ;
        RECT  2.255 0.705 2.310 0.875 ;
        RECT  2.195 1.515 2.310 1.945 ;
        RECT  1.160 1.515 2.195 1.655 ;
        RECT  0.990 1.515 1.160 1.945 ;
        END
        AntennaDiffArea 0.513 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.015 2.190 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.020 0.450 1.375 ;
        RECT  0.070 1.145 0.330 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.040 0.935 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.065 1.840 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.015 1.350 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.005 -0.210 2.520 0.210 ;
        RECT  0.835 -0.210 1.005 0.630 ;
        RECT  0.265 -0.210 0.835 0.210 ;
        RECT  0.095 -0.210 0.265 0.840 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.945 2.310 2.520 2.730 ;
        RECT  1.775 1.775 1.945 2.730 ;
        RECT  0.375 2.310 1.775 2.730 ;
        RECT  0.375 1.540 0.420 1.920 ;
        RECT  0.205 1.515 0.375 2.730 ;
        RECT  0.160 1.540 0.205 1.920 ;
        RECT  0.000 2.310 0.205 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  0.410 0.750 1.740 0.870 ;
    END
END OAI221X1AD
MACRO OAI221X2AD
    CLASS CORE ;
    FOREIGN OAI221X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.755 2.450 1.640 ;
        RECT  2.335 0.395 2.415 1.640 ;
        RECT  2.310 0.395 2.335 1.985 ;
        RECT  2.245 0.395 2.310 0.895 ;
        RECT  2.165 1.500 2.310 1.985 ;
        RECT  1.210 1.500 2.165 1.640 ;
        RECT  1.040 1.500 1.210 1.985 ;
        END
        AntennaDiffArea 0.839 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.880 1.015 2.190 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.145 0.470 1.375 ;
        RECT  0.320 1.030 0.440 1.375 ;
        RECT  0.070 1.145 0.320 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.015 0.800 1.935 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.015 1.760 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.015 1.350 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.040 -0.210 2.520 0.210 ;
        RECT  0.780 -0.210 1.040 0.390 ;
        RECT  0.255 -0.210 0.780 0.210 ;
        RECT  0.085 -0.210 0.255 0.795 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.935 2.310 2.520 2.730 ;
        RECT  1.765 1.760 1.935 2.730 ;
        RECT  0.375 2.310 1.765 2.730 ;
        RECT  0.205 1.615 0.375 2.730 ;
        RECT  0.000 2.310 0.205 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.885 0.395 2.055 0.870 ;
        RECT  1.120 0.750 1.885 0.870 ;
        RECT  1.525 0.435 1.695 0.630 ;
        RECT  0.615 0.510 1.525 0.630 ;
        RECT  0.445 0.365 0.615 0.795 ;
    END
END OAI221X2AD
MACRO OAI221X4AD
    CLASS CORE ;
    FOREIGN OAI221X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.270 0.750 4.410 1.640 ;
        RECT  3.670 0.750 4.270 0.880 ;
        RECT  4.265 1.520 4.270 1.640 ;
        RECT  4.095 1.520 4.265 1.980 ;
        RECT  3.525 1.520 4.095 1.640 ;
        RECT  3.355 1.520 3.525 1.950 ;
        RECT  1.900 1.520 3.355 1.640 ;
        RECT  1.730 1.520 1.900 1.950 ;
        RECT  0.325 1.520 1.730 1.640 ;
        RECT  0.155 1.520 0.325 1.950 ;
        END
        AntennaDiffArea 1.348 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 1.050 4.070 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.110 1.170 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.410 0.860 1.530 1.280 ;
        RECT  0.490 0.860 1.410 0.980 ;
        RECT  0.350 0.860 0.490 1.280 ;
        RECT  0.310 1.020 0.350 1.280 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.910 2.970 1.160 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.230 1.020 3.350 1.400 ;
        RECT  2.230 1.280 3.230 1.400 ;
        RECT  2.030 1.065 2.230 1.400 ;
        RECT  1.710 1.090 2.030 1.210 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.345 -0.210 4.480 0.210 ;
        RECT  1.175 -0.210 1.345 0.500 ;
        RECT  0.625 -0.210 1.175 0.210 ;
        RECT  0.455 -0.210 0.625 0.500 ;
        RECT  0.000 -0.210 0.455 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.895 2.310 4.480 2.730 ;
        RECT  3.725 1.775 3.895 2.730 ;
        RECT  2.795 2.310 3.725 2.730 ;
        RECT  2.625 1.775 2.795 2.730 ;
        RECT  1.030 2.310 2.625 2.730 ;
        RECT  0.860 1.775 1.030 2.730 ;
        RECT  0.000 2.310 0.860 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
        LAYER M1 ;
        RECT  3.525 0.380 4.310 0.500 ;
        RECT  3.355 0.380 3.525 0.810 ;
        RECT  2.065 0.380 3.355 0.500 ;
        RECT  1.750 0.620 3.210 0.740 ;
        RECT  1.895 0.330 2.065 0.500 ;
        RECT  1.490 0.360 1.750 0.740 ;
        RECT  1.030 0.620 1.490 0.740 ;
        RECT  0.770 0.360 1.030 0.740 ;
        RECT  0.230 0.620 0.770 0.740 ;
        RECT  0.110 0.395 0.230 0.915 ;
    END
END OAI221X4AD
MACRO OAI221XLAD
    CLASS CORE ;
    FOREIGN OAI221XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.725 2.450 1.685 ;
        RECT  2.255 0.725 2.310 0.895 ;
        RECT  0.885 1.515 2.310 1.685 ;
        END
        AntennaDiffArea 0.362 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.970 1.015 2.190 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.020 0.450 1.375 ;
        RECT  0.070 1.145 0.330 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.040 0.935 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.020 1.790 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.015 1.350 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 -0.210 2.520 0.210 ;
        RECT  0.790 -0.210 1.050 0.630 ;
        RECT  0.265 -0.210 0.790 0.210 ;
        RECT  0.095 -0.210 0.265 0.895 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.025 2.310 2.520 2.730 ;
        RECT  1.855 1.805 2.025 2.730 ;
        RECT  0.375 2.310 1.855 2.730 ;
        RECT  0.205 1.565 0.375 2.730 ;
        RECT  0.000 2.310 0.205 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  0.410 0.750 1.740 0.870 ;
    END
END OAI221XLAD
MACRO OAI222X1AD
    CLASS CORE ;
    FOREIGN OAI222X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.675 2.730 1.655 ;
        RECT  2.590 0.675 2.650 1.895 ;
        RECT  2.090 0.675 2.590 0.815 ;
        RECT  2.390 1.515 2.590 1.895 ;
        RECT  1.115 1.775 2.390 1.895 ;
        RECT  0.945 1.495 1.115 1.925 ;
        END
        AntennaDiffArea 0.472 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 1.035 2.095 1.655 ;
        RECT  1.750 1.425 1.925 1.655 ;
        END
        AntennaGateArea 0.0904 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.020 2.470 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 1.090 0.490 1.375 ;
        RECT  0.070 1.145 0.230 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 0.945 0.790 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.010 1.730 1.270 ;
        RECT  1.470 1.010 1.610 1.655 ;
        END
        AntennaGateArea 0.0904 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.020 1.350 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.955 -0.210 2.800 0.210 ;
        RECT  0.785 -0.210 0.955 0.385 ;
        RECT  0.265 -0.210 0.785 0.210 ;
        RECT  0.095 -0.210 0.265 0.825 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.900 2.310 2.800 2.730 ;
        RECT  1.730 2.015 1.900 2.730 ;
        RECT  0.365 2.310 1.730 2.730 ;
        RECT  0.195 1.520 0.365 2.730 ;
        RECT  0.000 2.310 0.195 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  0.410 0.700 1.650 0.820 ;
    END
END OAI222X1AD
MACRO OAI222X2AD
    CLASS CORE ;
    FOREIGN OAI222X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.925 0.635 2.990 1.715 ;
        RECT  2.850 0.635 2.925 1.990 ;
        RECT  2.295 0.635 2.850 0.775 ;
        RECT  2.755 1.515 2.850 1.990 ;
        RECT  1.195 1.515 2.755 1.715 ;
        RECT  0.910 1.515 1.195 1.945 ;
        END
        AntennaDiffArea 0.876 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.915 2.450 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.570 0.915 2.730 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.020 0.510 1.375 ;
        RECT  0.070 1.145 0.390 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.090 1.030 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 1.015 2.170 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.015 1.610 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.045 -0.210 3.080 0.210 ;
        RECT  0.875 -0.210 1.045 0.525 ;
        RECT  0.325 -0.210 0.875 0.210 ;
        RECT  0.155 -0.210 0.325 0.825 ;
        RECT  0.000 -0.210 0.155 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.265 2.310 3.080 2.730 ;
        RECT  1.835 1.995 2.265 2.730 ;
        RECT  0.445 2.310 1.835 2.730 ;
        RECT  0.275 1.540 0.445 2.730 ;
        RECT  0.000 2.310 0.275 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  2.135 0.380 2.940 0.500 ;
        RECT  1.965 0.380 2.135 0.825 ;
        RECT  1.190 0.380 1.965 0.500 ;
        RECT  0.685 0.655 1.765 0.825 ;
        RECT  0.515 0.395 0.685 0.825 ;
    END
END OAI222X2AD
MACRO OAI222X4AD
    CLASS CORE ;
    FOREIGN OAI222X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.880 0.790 4.970 1.590 ;
        RECT  4.830 0.790 4.880 1.950 ;
        RECT  4.660 0.790 4.830 0.910 ;
        RECT  4.710 1.450 4.830 1.950 ;
        RECT  3.470 1.450 4.710 1.590 ;
        RECT  4.540 0.620 4.660 0.910 ;
        RECT  3.645 0.620 4.540 0.740 ;
        RECT  3.300 1.450 3.470 1.970 ;
        RECT  1.880 1.450 3.300 1.590 ;
        RECT  1.710 1.450 1.880 1.950 ;
        RECT  0.315 1.450 1.710 1.590 ;
        RECT  0.145 1.450 0.315 1.980 ;
        END
        AntennaDiffArea 1.514 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.805 1.100 4.175 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.415 1.070 4.700 1.240 ;
        RECT  4.295 0.860 4.415 1.240 ;
        RECT  3.685 0.860 4.295 0.980 ;
        RECT  3.565 0.860 3.685 1.330 ;
        RECT  3.505 0.980 3.565 1.330 ;
        RECT  3.385 1.190 3.505 1.330 ;
        END
        AntennaGateArea 0.3249 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.655 1.120 1.175 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.435 1.020 1.525 1.280 ;
        RECT  1.315 0.860 1.435 1.280 ;
        RECT  0.535 0.860 1.315 0.980 ;
        RECT  0.415 0.860 0.535 1.330 ;
        RECT  0.295 1.085 0.415 1.330 ;
        END
        AntennaGateArea 0.3249 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.420 1.100 2.940 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.145 0.860 3.265 1.280 ;
        RECT  2.185 0.860 3.145 0.980 ;
        RECT  1.805 0.860 2.185 1.260 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.340 -0.210 5.040 0.210 ;
        RECT  1.170 -0.210 1.340 0.465 ;
        RECT  0.615 -0.210 1.170 0.210 ;
        RECT  0.445 -0.210 0.615 0.465 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.220 2.310 5.040 2.730 ;
        RECT  4.050 1.735 4.220 2.730 ;
        RECT  2.760 2.310 4.050 2.730 ;
        RECT  2.590 1.735 2.760 2.730 ;
        RECT  0.975 2.310 2.590 2.730 ;
        RECT  0.805 1.735 0.975 2.730 ;
        RECT  0.000 2.310 0.805 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.040 2.520 ;
        LAYER M1 ;
        RECT  4.795 0.380 4.915 0.640 ;
        RECT  2.060 0.380 4.795 0.500 ;
        RECT  1.745 0.620 3.185 0.740 ;
        RECT  1.890 0.330 2.060 0.500 ;
        RECT  1.485 0.360 1.745 0.740 ;
        RECT  1.020 0.620 1.485 0.740 ;
        RECT  0.760 0.360 1.020 0.740 ;
        RECT  0.255 0.620 0.760 0.740 ;
        RECT  0.085 0.410 0.255 0.840 ;
    END
END OAI222X4AD
MACRO OAI222XLAD
    CLASS CORE ;
    FOREIGN OAI222XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.605 0.740 2.730 1.655 ;
        RECT  2.590 0.740 2.605 1.685 ;
        RECT  2.090 0.740 2.590 0.880 ;
        RECT  2.555 1.515 2.590 1.685 ;
        RECT  2.435 1.515 2.555 1.895 ;
        RECT  1.115 1.775 2.435 1.895 ;
        RECT  0.995 1.495 1.115 1.895 ;
        RECT  0.945 1.495 0.995 1.665 ;
        END
        AntennaDiffArea 0.312 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.925 1.020 2.095 1.655 ;
        RECT  1.750 1.425 1.925 1.655 ;
        END
        AntennaGateArea 0.0602 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.020 2.470 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.230 1.090 0.490 1.375 ;
        RECT  0.070 1.145 0.230 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.010 0.790 1.440 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.010 1.730 1.270 ;
        RECT  1.470 1.010 1.610 1.655 ;
        END
        AntennaGateArea 0.0602 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.020 1.350 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.955 -0.210 2.800 0.210 ;
        RECT  0.785 -0.210 0.955 0.475 ;
        RECT  0.265 -0.210 0.785 0.210 ;
        RECT  0.095 -0.210 0.265 0.905 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.900 2.310 2.800 2.730 ;
        RECT  1.730 2.015 1.900 2.730 ;
        RECT  0.355 2.310 1.730 2.730 ;
        RECT  0.185 1.495 0.355 2.730 ;
        RECT  0.000 2.310 0.185 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  0.410 0.760 1.650 0.880 ;
    END
END OAI222XLAD
MACRO OAI22X1AD
    CLASS CORE ;
    FOREIGN OAI22X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.640 1.295 1.000 ;
        RECT  0.490 0.880 1.125 1.000 ;
        RECT  0.490 1.730 0.980 1.935 ;
        RECT  0.370 0.880 0.490 1.935 ;
        RECT  0.350 1.705 0.370 1.935 ;
        END
        AntennaDiffArea 0.234 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.070 0.230 1.530 ;
        END
        AntennaGateArea 0.09 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.615 1.120 0.785 1.540 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.640 1.610 1.315 ;
        RECT  1.255 1.145 1.470 1.315 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.090 1.470 1.375 1.610 ;
        RECT  0.915 1.120 1.090 1.610 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.555 -0.210 1.680 0.210 ;
        RECT  0.385 -0.210 0.555 0.360 ;
        RECT  0.000 -0.210 0.385 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.545 2.310 1.680 2.730 ;
        RECT  1.375 1.780 1.545 2.730 ;
        RECT  0.230 2.310 1.375 2.730 ;
        RECT  0.110 1.670 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  0.255 0.640 0.980 0.760 ;
        RECT  0.085 0.640 0.255 0.810 ;
    END
END OAI22X1AD
MACRO OAI22X2AD
    CLASS CORE ;
    FOREIGN OAI22X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.325 0.665 1.510 0.900 ;
        RECT  0.640 0.780 1.325 0.900 ;
        RECT  0.965 1.495 1.135 1.955 ;
        RECT  0.640 1.495 0.965 1.695 ;
        RECT  0.520 0.780 0.640 1.695 ;
        RECT  0.350 0.780 0.520 1.095 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.020 0.230 1.490 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.760 1.020 1.050 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.040 1.890 1.375 ;
        RECT  1.505 1.040 1.750 1.300 ;
        END
        AntennaGateArea 0.1629 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.020 1.385 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.700 -0.210 1.960 0.210 ;
        RECT  0.530 -0.210 0.700 0.415 ;
        RECT  0.000 -0.210 0.530 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.795 2.310 1.960 2.730 ;
        RECT  1.625 1.585 1.795 2.730 ;
        RECT  0.400 2.310 1.625 2.730 ;
        RECT  0.230 1.635 0.400 2.730 ;
        RECT  0.000 2.310 0.230 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.695 0.395 1.865 0.840 ;
        RECT  1.145 0.395 1.695 0.515 ;
        RECT  0.960 0.395 1.145 0.660 ;
        RECT  0.230 0.540 0.960 0.660 ;
        RECT  0.110 0.370 0.230 0.890 ;
    END
END OAI22X2AD
MACRO OAI22X4AD
    CLASS CORE ;
    FOREIGN OAI22X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.835 3.290 1.820 ;
        RECT  2.845 0.835 3.150 0.965 ;
        RECT  2.485 1.690 3.150 1.820 ;
        RECT  2.675 0.630 2.845 0.965 ;
        RECT  2.125 0.835 2.675 0.965 ;
        RECT  2.315 1.690 2.485 2.140 ;
        RECT  0.985 1.690 2.315 1.820 ;
        RECT  1.955 0.630 2.125 0.965 ;
        RECT  0.815 1.690 0.985 2.135 ;
        END
        AntennaDiffArea 0.85 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.420 1.110 1.570 1.230 ;
        RECT  1.280 1.110 1.420 1.570 ;
        RECT  0.490 1.450 1.280 1.570 ;
        RECT  0.220 1.110 0.490 1.655 ;
        END
        AntennaGateArea 0.3249 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.110 1.150 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 1.085 3.010 1.570 ;
        RECT  1.990 1.450 2.835 1.570 ;
        RECT  1.730 1.090 1.990 1.570 ;
        END
        AntennaGateArea 0.3249 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 1.090 2.650 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.365 -0.210 3.360 0.210 ;
        RECT  1.195 -0.210 1.365 0.690 ;
        RECT  0.625 -0.210 1.195 0.210 ;
        RECT  0.455 -0.210 0.625 0.680 ;
        RECT  0.000 -0.210 0.455 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.145 2.310 3.360 2.730 ;
        RECT  2.975 1.970 3.145 2.730 ;
        RECT  1.745 2.310 2.975 2.730 ;
        RECT  1.575 1.995 1.745 2.730 ;
        RECT  0.325 2.310 1.575 2.730 ;
        RECT  0.155 1.775 0.325 2.730 ;
        RECT  0.000 2.310 0.155 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  3.045 0.380 3.215 0.665 ;
        RECT  2.485 0.380 3.045 0.510 ;
        RECT  2.315 0.380 2.485 0.615 ;
        RECT  1.765 0.380 2.315 0.510 ;
        RECT  1.595 0.380 1.765 0.955 ;
        RECT  0.985 0.835 1.595 0.955 ;
        RECT  0.815 0.435 0.985 0.955 ;
        RECT  0.255 0.835 0.815 0.955 ;
        RECT  0.085 0.410 0.255 0.955 ;
    END
END OAI22X4AD
MACRO OAI22XLAD
    CLASS CORE ;
    FOREIGN OAI22XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.125 0.640 1.295 1.025 ;
        RECT  0.490 0.905 1.125 1.025 ;
        RECT  0.490 1.730 0.980 1.935 ;
        RECT  0.350 0.905 0.490 1.935 ;
        END
        AntennaDiffArea 0.156 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.145 0.230 1.530 ;
        END
        AntennaGateArea 0.06 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.615 1.145 0.785 1.540 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.640 1.610 1.315 ;
        RECT  1.255 1.145 1.470 1.315 ;
        END
        AntennaGateArea 0.06 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.090 1.470 1.375 1.610 ;
        RECT  0.915 1.145 1.090 1.610 ;
        END
        AntennaGateArea 0.06 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.555 -0.210 1.680 0.210 ;
        RECT  0.385 -0.210 0.555 0.380 ;
        RECT  0.000 -0.210 0.385 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.595 2.310 1.680 2.730 ;
        RECT  1.425 1.730 1.595 2.730 ;
        RECT  0.230 2.310 1.425 2.730 ;
        RECT  0.110 1.650 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  0.255 0.665 0.980 0.785 ;
        RECT  0.085 0.640 0.255 0.810 ;
    END
END OAI22XLAD
MACRO OAI2B11X1AD
    CLASS CORE ;
    FOREIGN OAI2B11X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.155 0.670 2.170 1.375 ;
        RECT  2.010 0.670 2.155 1.925 ;
        RECT  1.985 1.495 2.010 1.925 ;
        RECT  1.435 1.495 1.985 1.615 ;
        RECT  1.265 1.495 1.435 1.925 ;
        END
        AntennaDiffArea 0.365 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.865 1.690 1.285 ;
        END
        AntennaGateArea 0.09 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.705 0.350 2.135 0.510 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.335 1.025 0.550 1.375 ;
        END
        AntennaGateArea 0.041 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.035 1.320 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.185 -0.210 2.240 0.210 ;
        RECT  1.015 -0.210 1.185 0.845 ;
        RECT  0.555 -0.210 1.015 0.210 ;
        RECT  0.385 -0.210 0.555 0.470 ;
        RECT  0.000 -0.210 0.385 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.795 2.310 2.240 2.730 ;
        RECT  1.625 1.750 1.795 2.730 ;
        RECT  0.775 2.310 1.625 2.730 ;
        RECT  0.605 1.525 0.775 2.730 ;
        RECT  0.000 2.310 0.605 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  0.670 0.785 0.790 1.285 ;
        RECT  0.265 0.785 0.670 0.905 ;
        RECT  0.215 1.490 0.285 1.660 ;
        RECT  0.215 0.735 0.265 0.905 ;
        RECT  0.095 0.735 0.215 1.660 ;
    END
END OAI2B11X1AD
MACRO OAI2B11X2AD
    CLASS CORE ;
    FOREIGN OAI2B11X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.975 0.355 2.145 0.785 ;
        RECT  1.975 1.515 2.145 1.990 ;
        RECT  1.890 0.585 1.975 0.785 ;
        RECT  1.890 1.515 1.975 1.635 ;
        RECT  1.750 0.585 1.890 1.635 ;
        RECT  1.425 1.515 1.750 1.635 ;
        RECT  1.255 1.515 1.425 1.990 ;
        END
        AntennaDiffArea 0.615 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.410 1.015 1.610 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.935 2.170 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.285 1.705 0.490 2.050 ;
        END
        AntennaGateArea 0.0653 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.015 1.260 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.220 -0.210 2.240 0.210 ;
        RECT  0.960 -0.210 1.220 0.650 ;
        RECT  0.255 -0.210 0.960 0.210 ;
        RECT  0.085 -0.210 0.255 0.405 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.785 2.310 2.240 2.730 ;
        RECT  1.615 1.780 1.785 2.730 ;
        RECT  0.740 2.310 1.615 2.730 ;
        RECT  0.620 1.640 0.740 2.730 ;
        RECT  0.000 2.310 0.620 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.365 0.375 1.535 0.890 ;
        RECT  0.815 0.770 1.365 0.890 ;
        RECT  0.695 0.340 0.815 0.890 ;
        RECT  0.520 1.020 0.790 1.280 ;
        RECT  0.645 0.340 0.695 0.510 ;
        RECT  0.400 0.690 0.520 1.495 ;
        RECT  0.365 1.375 0.400 1.495 ;
        RECT  0.195 1.375 0.365 1.545 ;
    END
END OAI2B11X2AD
MACRO OAI2B11X4AD
    CLASS CORE ;
    FOREIGN OAI2B11X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.825 0.665 3.850 1.655 ;
        RECT  3.710 0.665 3.825 1.975 ;
        RECT  2.890 0.665 3.710 0.785 ;
        RECT  3.655 1.525 3.710 1.975 ;
        RECT  3.105 1.525 3.655 1.655 ;
        RECT  2.935 1.525 3.105 1.975 ;
        RECT  2.320 1.525 2.935 1.655 ;
        RECT  2.150 1.525 2.320 1.975 ;
        RECT  1.030 1.525 2.150 1.655 ;
        RECT  0.860 1.525 1.030 2.020 ;
        END
        AntennaDiffArea 1.092 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.470 1.015 3.590 1.405 ;
        RECT  2.570 1.285 3.470 1.405 ;
        RECT  2.265 1.020 2.570 1.405 ;
        END
        AntennaGateArea 0.324 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 0.905 3.210 1.165 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.015 0.375 1.230 ;
        RECT  0.070 1.015 0.210 1.375 ;
        END
        AntennaGateArea 0.129 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.025 0.880 2.145 1.275 ;
        RECT  1.195 0.880 2.025 1.000 ;
        RECT  0.865 0.880 1.195 1.165 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.070 -0.210 3.920 0.210 ;
        RECT  1.900 -0.210 2.070 0.480 ;
        RECT  1.350 -0.210 1.900 0.210 ;
        RECT  1.180 -0.210 1.350 0.480 ;
        RECT  0.255 -0.210 1.180 0.210 ;
        RECT  0.085 -0.210 0.255 0.845 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.465 2.310 3.920 2.730 ;
        RECT  3.295 1.845 3.465 2.730 ;
        RECT  2.690 2.310 3.295 2.730 ;
        RECT  2.520 1.845 2.690 2.730 ;
        RECT  1.710 2.310 2.520 2.730 ;
        RECT  1.540 1.845 1.710 2.730 ;
        RECT  0.255 2.310 1.540 2.730 ;
        RECT  0.085 1.505 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  2.430 0.425 3.810 0.545 ;
        RECT  2.260 0.330 2.430 0.760 ;
        RECT  1.710 0.640 2.260 0.760 ;
        RECT  1.435 1.120 1.875 1.240 ;
        RECT  1.540 0.330 1.710 0.760 ;
        RECT  0.990 0.640 1.540 0.760 ;
        RECT  1.315 1.120 1.435 1.405 ;
        RECT  0.615 1.285 1.315 1.405 ;
        RECT  0.820 0.330 0.990 0.760 ;
        RECT  0.495 0.415 0.615 1.920 ;
        RECT  0.445 0.415 0.495 0.845 ;
        RECT  0.445 1.490 0.495 1.920 ;
    END
END OAI2B11X4AD
MACRO OAI2B11XLAD
    CLASS CORE ;
    FOREIGN OAI2B11XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.685 2.170 1.375 ;
        RECT  2.010 0.685 2.130 1.820 ;
        RECT  1.435 1.495 2.010 1.615 ;
        RECT  1.315 1.495 1.435 1.775 ;
        RECT  1.265 1.605 1.315 1.775 ;
        END
        AntennaDiffArea 0.242 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.865 1.690 1.285 ;
        END
        AntennaGateArea 0.06 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.705 0.350 2.135 0.565 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.335 1.025 0.550 1.375 ;
        END
        AntennaGateArea 0.04 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.035 1.320 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.185 -0.210 2.240 0.210 ;
        RECT  1.015 -0.210 1.185 0.900 ;
        RECT  0.545 -0.210 1.015 0.210 ;
        RECT  0.375 -0.210 0.545 0.470 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.840 2.310 2.240 2.730 ;
        RECT  1.580 1.735 1.840 2.730 ;
        RECT  0.755 2.310 1.580 2.730 ;
        RECT  0.585 1.525 0.755 2.730 ;
        RECT  0.000 2.310 0.585 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  0.670 0.785 0.790 1.285 ;
        RECT  0.265 0.785 0.670 0.905 ;
        RECT  0.215 1.510 0.285 1.680 ;
        RECT  0.215 0.735 0.265 0.905 ;
        RECT  0.095 0.735 0.215 1.680 ;
    END
END OAI2B11XLAD
MACRO OAI2B1X1AD
    CLASS CORE ;
    FOREIGN OAI2B1X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.770 0.585 1.890 1.895 ;
        RECT  1.720 0.585 1.770 0.890 ;
        RECT  1.460 1.775 1.770 1.895 ;
        RECT  1.200 1.775 1.460 2.155 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.455 1.245 1.650 1.655 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.345 0.710 0.495 1.230 ;
        END
        AntennaGateArea 0.0415 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 1.240 1.330 1.655 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.175 -0.210 1.960 0.210 ;
        RECT  0.485 -0.210 1.175 0.385 ;
        RECT  0.000 -0.210 0.485 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.775 2.310 1.960 2.730 ;
        RECT  1.605 2.015 1.775 2.730 ;
        RECT  0.735 2.310 1.605 2.730 ;
        RECT  0.565 1.655 0.735 2.730 ;
        RECT  0.000 2.310 0.565 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.455 0.735 1.505 0.905 ;
        RECT  1.335 0.735 1.455 1.120 ;
        RECT  0.840 1.000 1.335 1.120 ;
        RECT  0.275 1.350 0.950 1.470 ;
        RECT  0.720 0.735 0.840 1.120 ;
        RECT  0.645 0.735 0.720 0.905 ;
        RECT  0.225 0.350 0.275 0.520 ;
        RECT  0.225 1.350 0.275 1.775 ;
        RECT  0.105 0.350 0.225 1.775 ;
    END
END OAI2B1X1AD
MACRO OAI2B1X2AD
    CLASS CORE ;
    FOREIGN OAI2B1X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.865 2.170 1.375 ;
        RECT  2.010 0.405 2.130 1.625 ;
        RECT  1.960 0.405 2.010 0.835 ;
        RECT  1.700 1.505 2.010 1.625 ;
        RECT  1.530 1.505 1.700 2.015 ;
        END
        AntennaDiffArea 0.401 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 1.015 1.890 1.375 ;
        END
        AntennaGateArea 0.1629 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.255 1.020 0.375 1.375 ;
        RECT  0.070 1.115 0.255 1.375 ;
        END
        AntennaGateArea 0.0654 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.065 1.530 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.450 -0.210 2.240 0.210 ;
        RECT  1.190 -0.210 1.450 0.650 ;
        RECT  0.330 -0.210 1.190 0.210 ;
        RECT  0.160 -0.210 0.330 0.865 ;
        RECT  0.000 -0.210 0.160 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.060 2.310 2.240 2.730 ;
        RECT  1.890 1.790 2.060 2.730 ;
        RECT  1.040 2.310 1.890 2.730 ;
        RECT  0.870 1.635 1.040 2.730 ;
        RECT  0.000 2.310 0.870 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.600 0.405 1.770 0.895 ;
        RECT  1.040 0.775 1.600 0.895 ;
        RECT  0.640 1.065 1.070 1.235 ;
        RECT  0.870 0.410 1.040 0.895 ;
        RECT  0.640 0.695 0.690 0.865 ;
        RECT  0.520 0.695 0.640 1.675 ;
        RECT  0.330 1.555 0.520 1.675 ;
        RECT  0.160 1.555 0.330 1.725 ;
    END
END OAI2B1X2AD
MACRO OAI2B1X4AD
    CLASS CORE ;
    FOREIGN OAI2B1X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.725 3.290 1.580 ;
        RECT  2.880 0.725 3.150 0.855 ;
        RECT  2.880 1.450 3.150 1.580 ;
        RECT  2.710 0.685 2.880 0.855 ;
        RECT  2.710 1.450 2.880 2.035 ;
        RECT  1.800 1.450 2.710 1.580 ;
        RECT  1.630 1.450 1.800 2.000 ;
        END
        AntennaDiffArea 0.664 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.510 1.080 2.870 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.980 0.440 1.375 ;
        RECT  0.070 1.145 0.320 1.375 ;
        END
        AntennaGateArea 0.129 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 1.120 1.965 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.160 -0.210 3.360 0.210 ;
        RECT  1.990 -0.210 2.160 0.510 ;
        RECT  1.440 -0.210 1.990 0.210 ;
        RECT  1.270 -0.210 1.440 0.510 ;
        RECT  0.370 -0.210 1.270 0.210 ;
        RECT  0.200 -0.210 0.370 0.860 ;
        RECT  0.000 -0.210 0.200 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.240 2.310 3.360 2.730 ;
        RECT  3.070 1.725 3.240 2.730 ;
        RECT  2.490 2.310 3.070 2.730 ;
        RECT  2.320 1.725 2.490 2.730 ;
        RECT  1.065 2.310 2.320 2.730 ;
        RECT  0.875 1.605 1.065 2.730 ;
        RECT  0.000 2.310 0.875 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  3.070 0.380 3.240 0.550 ;
        RECT  2.520 0.380 3.070 0.500 ;
        RECT  2.350 0.330 2.520 0.760 ;
        RECT  2.215 1.090 2.355 1.210 ;
        RECT  1.800 0.640 2.350 0.760 ;
        RECT  2.095 0.880 2.215 1.210 ;
        RECT  1.260 0.880 2.095 1.000 ;
        RECT  1.630 0.330 1.800 0.760 ;
        RECT  1.080 0.640 1.630 0.760 ;
        RECT  1.090 0.880 1.260 1.235 ;
        RECT  0.730 1.065 1.090 1.235 ;
        RECT  0.910 0.330 1.080 0.760 ;
        RECT  0.560 0.435 0.730 1.615 ;
        RECT  0.370 1.495 0.560 1.615 ;
        RECT  0.200 1.495 0.370 2.010 ;
    END
END OAI2B1X4AD
MACRO OAI2B1XLAD
    CLASS CORE ;
    FOREIGN OAI2B1XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.770 0.690 1.890 1.895 ;
        RECT  1.720 0.690 1.770 1.095 ;
        RECT  1.415 1.775 1.770 1.895 ;
        RECT  1.245 1.775 1.415 1.945 ;
        END
        AntennaDiffArea 0.15 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.455 1.245 1.650 1.655 ;
        END
        AntennaGateArea 0.0604 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.345 0.685 0.495 1.205 ;
        END
        AntennaGateArea 0.04 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 1.240 1.330 1.655 ;
        END
        AntennaGateArea 0.06 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.165 -0.210 1.960 0.210 ;
        RECT  0.995 -0.210 1.165 0.475 ;
        RECT  0.655 -0.210 0.995 0.210 ;
        RECT  0.485 -0.210 0.655 0.565 ;
        RECT  0.000 -0.210 0.485 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.840 2.310 1.960 2.730 ;
        RECT  1.580 2.015 1.840 2.730 ;
        RECT  0.715 2.310 1.580 2.730 ;
        RECT  0.545 1.595 0.715 2.730 ;
        RECT  0.000 2.310 0.545 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.455 0.735 1.505 0.905 ;
        RECT  1.335 0.735 1.455 1.120 ;
        RECT  0.810 1.000 1.335 1.120 ;
        RECT  0.275 1.325 0.950 1.445 ;
        RECT  0.690 0.735 0.810 1.120 ;
        RECT  0.615 0.735 0.690 0.905 ;
        RECT  0.225 0.395 0.275 0.565 ;
        RECT  0.225 1.325 0.275 1.765 ;
        RECT  0.105 0.395 0.225 1.765 ;
    END
END OAI2B1XLAD
MACRO OAI2B2X1AD
    CLASS CORE ;
    FOREIGN OAI2B2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.210 0.585 1.330 1.615 ;
        RECT  1.140 0.585 1.210 0.855 ;
        RECT  0.905 1.495 1.210 1.615 ;
        RECT  1.045 0.685 1.140 0.855 ;
        RECT  0.735 1.495 0.905 1.955 ;
        END
        AntennaDiffArea 0.234 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.245 1.050 0.415 1.220 ;
        RECT  0.210 1.100 0.245 1.220 ;
        RECT  0.070 1.100 0.210 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.000 0.770 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.025 1.900 1.375 ;
        END
        AntennaGateArea 0.041 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.000 1.085 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.845 -0.210 2.240 0.210 ;
        RECT  1.675 -0.210 1.845 0.475 ;
        RECT  0.545 -0.210 1.675 0.210 ;
        RECT  0.375 -0.210 0.545 0.855 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.620 2.310 2.240 2.730 ;
        RECT  1.450 1.495 1.620 2.730 ;
        RECT  0.295 2.310 1.450 2.730 ;
        RECT  0.125 1.525 0.295 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  2.020 0.735 2.140 1.615 ;
        RECT  1.965 0.735 2.020 0.905 ;
        RECT  1.860 1.495 2.020 1.615 ;
        RECT  1.570 0.735 1.965 0.855 ;
        RECT  1.450 0.735 1.570 1.265 ;
    END
END OAI2B2X1AD
MACRO OAI2B2X2AD
    CLASS CORE ;
    FOREIGN OAI2B2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.255 0.630 1.375 1.895 ;
        RECT  1.145 0.630 1.255 0.850 ;
        RECT  1.050 1.775 1.255 1.895 ;
        RECT  0.790 1.775 1.050 2.155 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.260 1.025 0.435 1.195 ;
        RECT  0.210 1.075 0.260 1.195 ;
        RECT  0.070 1.075 0.210 1.655 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.010 0.770 1.655 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.215 1.145 2.450 1.375 ;
        RECT  1.835 1.020 2.215 1.375 ;
        END
        AntennaGateArea 0.065 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.010 1.070 1.655 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.415 -0.210 2.520 0.210 ;
        RECT  2.245 -0.210 2.415 0.835 ;
        RECT  0.690 -0.210 2.245 0.210 ;
        RECT  0.430 -0.210 0.690 0.650 ;
        RECT  0.000 -0.210 0.430 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.665 2.310 2.520 2.730 ;
        RECT  1.495 1.755 1.665 2.730 ;
        RECT  0.345 2.310 1.495 2.730 ;
        RECT  0.175 1.780 0.345 2.730 ;
        RECT  0.000 2.310 0.175 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.960 1.495 2.130 1.665 ;
        RECT  1.885 0.725 2.055 0.895 ;
        RECT  1.615 1.495 1.960 1.615 ;
        RECT  1.615 0.775 1.885 0.895 ;
        RECT  1.555 0.340 1.725 0.510 ;
        RECT  1.495 0.775 1.615 1.615 ;
        RECT  1.005 0.390 1.555 0.510 ;
        RECT  0.835 0.390 1.005 0.890 ;
        RECT  0.285 0.770 0.835 0.890 ;
        RECT  0.115 0.410 0.285 0.890 ;
    END
END OAI2B2X2AD
MACRO OAI2B2X4AD
    CLASS CORE ;
    FOREIGN OAI2B2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.635 0.670 2.805 0.840 ;
        RECT  2.085 0.670 2.635 0.800 ;
        RECT  2.275 1.710 2.445 2.140 ;
        RECT  1.665 1.750 2.275 1.890 ;
        RECT  2.035 0.670 2.085 0.840 ;
        RECT  1.915 0.670 2.035 0.965 ;
        RECT  1.665 0.845 1.915 0.965 ;
        RECT  1.545 0.845 1.665 1.890 ;
        RECT  1.000 1.750 1.545 1.890 ;
        RECT  0.830 1.705 1.000 2.135 ;
        END
        AntennaDiffArea 0.844 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.305 0.995 1.425 1.570 ;
        RECT  0.490 1.450 1.305 1.570 ;
        RECT  0.320 1.110 0.490 1.570 ;
        RECT  0.230 1.110 0.320 1.230 ;
        END
        AntennaGateArea 0.324 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.645 1.110 1.165 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.105 1.065 3.365 1.330 ;
        END
        AntennaGateArea 0.1294 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.585 1.090 2.670 1.210 ;
        RECT  2.150 1.090 2.585 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.475 -0.210 3.920 0.210 ;
        RECT  3.305 -0.210 3.475 0.905 ;
        RECT  1.365 -0.210 3.305 0.210 ;
        RECT  1.195 -0.210 1.365 0.470 ;
        RECT  0.640 -0.210 1.195 0.210 ;
        RECT  0.470 -0.210 0.640 0.675 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.105 2.310 3.920 2.730 ;
        RECT  2.935 1.690 3.105 2.730 ;
        RECT  1.715 2.310 2.935 2.730 ;
        RECT  1.545 2.045 1.715 2.730 ;
        RECT  0.340 2.310 1.545 2.730 ;
        RECT  0.170 1.735 0.340 2.730 ;
        RECT  0.000 2.310 0.170 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  3.785 0.440 3.835 0.870 ;
        RECT  3.665 0.440 3.785 1.570 ;
        RECT  3.485 1.450 3.665 1.570 ;
        RECT  3.315 1.450 3.485 1.880 ;
        RECT  2.930 1.450 3.315 1.570 ;
        RECT  2.995 0.390 3.165 0.560 ;
        RECT  1.725 0.390 2.995 0.520 ;
        RECT  2.810 1.020 2.930 1.570 ;
        RECT  1.965 1.450 2.810 1.570 ;
        RECT  1.845 1.085 1.965 1.570 ;
        RECT  1.795 1.085 1.845 1.255 ;
        RECT  1.555 0.390 1.725 0.720 ;
        RECT  1.000 0.600 1.555 0.720 ;
        RECT  0.830 0.435 1.000 0.955 ;
        RECT  0.280 0.835 0.830 0.955 ;
        RECT  0.110 0.410 0.280 0.955 ;
    END
END OAI2B2X4AD
MACRO OAI2B2XLAD
    CLASS CORE ;
    FOREIGN OAI2B2XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.210 0.585 1.330 1.895 ;
        RECT  0.910 0.585 1.210 0.840 ;
        RECT  0.905 1.775 1.210 1.895 ;
        RECT  0.735 1.775 0.905 1.945 ;
        END
        AntennaDiffArea 0.156 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 0.960 0.420 1.480 ;
        RECT  0.070 1.145 0.300 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 0.960 0.770 1.655 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.025 1.900 1.375 ;
        END
        AntennaGateArea 0.04 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.960 1.085 1.655 ;
        END
        AntennaGateArea 0.06 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.845 -0.210 2.240 0.210 ;
        RECT  1.675 -0.210 1.845 0.475 ;
        RECT  0.590 -0.210 1.675 0.210 ;
        RECT  0.330 -0.210 0.590 0.840 ;
        RECT  0.000 -0.210 0.330 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.620 2.310 2.240 2.730 ;
        RECT  1.450 1.575 1.620 2.730 ;
        RECT  0.295 2.310 1.450 2.730 ;
        RECT  0.125 1.775 0.295 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  2.020 0.735 2.140 1.745 ;
        RECT  1.965 0.735 2.020 0.905 ;
        RECT  1.905 1.575 2.020 1.745 ;
        RECT  1.570 0.735 1.965 0.855 ;
        RECT  1.450 0.735 1.570 1.265 ;
    END
END OAI2B2XLAD
MACRO OAI2BB1X1AD
    CLASS CORE ;
    FOREIGN OAI2BB1X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.490 0.640 1.610 1.655 ;
        RECT  1.430 0.640 1.490 0.900 ;
        RECT  1.460 1.425 1.490 1.655 ;
        RECT  1.225 1.525 1.460 1.655 ;
        RECT  1.055 1.525 1.225 1.955 ;
        END
        AntennaDiffArea 0.235 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.020 1.070 1.405 ;
        END
        AntennaGateArea 0.091 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.250 1.280 ;
        RECT  0.070 1.020 0.210 1.630 ;
        END
        AntennaGateArea 0.0433 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.020 0.790 1.375 ;
        END
        AntennaGateArea 0.0434 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.905 -0.210 1.680 0.210 ;
        RECT  0.735 -0.210 0.905 0.660 ;
        RECT  0.000 -0.210 0.735 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.585 2.310 1.680 2.730 ;
        RECT  1.415 1.815 1.585 2.730 ;
        RECT  0.805 2.310 1.415 2.730 ;
        RECT  0.115 1.905 0.805 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.310 1.020 1.370 1.280 ;
        RECT  1.190 0.780 1.310 1.280 ;
        RECT  0.490 0.780 1.190 0.900 ;
        RECT  0.490 1.500 0.600 1.620 ;
        RECT  0.370 0.780 0.490 1.620 ;
        RECT  0.265 0.780 0.370 0.900 ;
        RECT  0.340 1.500 0.370 1.620 ;
        RECT  0.095 0.730 0.265 0.900 ;
    END
END OAI2BB1X1AD
MACRO OAI2BB1X2AD
    CLASS CORE ;
    FOREIGN OAI2BB1X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.860 1.145 1.890 1.375 ;
        RECT  1.795 0.640 1.860 1.555 ;
        RECT  1.740 0.430 1.795 1.555 ;
        RECT  1.625 0.430 1.740 0.860 ;
        RECT  1.495 1.435 1.740 1.555 ;
        RECT  1.325 1.435 1.495 1.985 ;
        END
        AntennaDiffArea 0.401 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 1.020 1.265 1.280 ;
        RECT  0.910 1.020 1.115 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.020 0.270 1.385 ;
        RECT  0.070 1.145 0.130 1.385 ;
        END
        AntennaGateArea 0.0774 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.970 0.790 1.375 ;
        END
        AntennaGateArea 0.077 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.180 -0.210 1.960 0.210 ;
        RECT  0.750 -0.210 1.180 0.610 ;
        RECT  0.000 -0.210 0.750 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.855 2.310 1.960 2.730 ;
        RECT  1.685 1.725 1.855 2.730 ;
        RECT  1.135 2.310 1.685 2.730 ;
        RECT  0.965 1.625 1.135 2.730 ;
        RECT  0.270 2.310 0.965 2.730 ;
        RECT  0.100 1.505 0.270 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.505 1.000 1.620 1.260 ;
        RECT  1.385 0.730 1.505 1.260 ;
        RECT  0.510 0.730 1.385 0.850 ;
        RECT  0.510 1.495 0.650 1.665 ;
        RECT  0.390 0.730 0.510 1.665 ;
        RECT  0.290 0.730 0.390 0.850 ;
        RECT  0.120 0.680 0.290 0.850 ;
    END
END OAI2BB1X2AD
MACRO OAI2BB1X4AD
    CLASS CORE ;
    FOREIGN OAI2BB1X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.410 1.005 2.450 1.515 ;
        RECT  2.280 0.770 2.410 1.695 ;
        RECT  1.695 0.770 2.280 0.900 ;
        RECT  2.055 1.565 2.280 1.695 ;
        RECT  1.885 1.565 2.055 1.995 ;
        RECT  1.335 1.565 1.885 1.695 ;
        RECT  1.525 0.430 1.695 0.900 ;
        RECT  1.165 1.565 1.335 1.995 ;
        END
        AntennaDiffArea 0.664 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.020 2.150 1.435 ;
        RECT  1.160 1.315 2.030 1.435 ;
        RECT  1.040 1.020 1.160 1.435 ;
        RECT  0.910 1.020 1.040 1.410 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.260 1.280 ;
        RECT  0.130 1.020 0.210 1.420 ;
        RECT  0.070 1.145 0.130 1.420 ;
        END
        AntennaGateArea 0.147 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.020 0.790 1.420 ;
        END
        AntennaGateArea 0.147 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.410 -0.210 2.520 0.210 ;
        RECT  2.150 -0.210 2.410 0.650 ;
        RECT  1.015 -0.210 2.150 0.210 ;
        RECT  0.755 -0.210 1.015 0.650 ;
        RECT  0.000 -0.210 0.755 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.415 2.310 2.520 2.730 ;
        RECT  2.245 1.855 2.415 2.730 ;
        RECT  1.695 2.310 2.245 2.730 ;
        RECT  1.525 1.865 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.575 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.540 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.495 1.050 1.880 1.170 ;
        RECT  1.400 1.025 1.495 1.170 ;
        RECT  1.360 0.780 1.400 1.170 ;
        RECT  1.280 0.780 1.360 1.145 ;
        RECT  0.500 0.780 1.280 0.900 ;
        RECT  0.500 1.540 0.615 1.970 ;
        RECT  0.380 0.780 0.500 1.970 ;
        RECT  0.255 0.780 0.380 0.900 ;
        RECT  0.085 0.445 0.255 0.900 ;
    END
END OAI2BB1X4AD
MACRO OAI2BB1XLAD
    CLASS CORE ;
    FOREIGN OAI2BB1XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.490 0.685 1.610 1.655 ;
        RECT  1.430 0.685 1.490 0.945 ;
        RECT  1.460 1.425 1.490 1.655 ;
        RECT  1.225 1.535 1.460 1.655 ;
        RECT  1.055 1.535 1.225 1.825 ;
        END
        AntennaDiffArea 0.157 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.020 1.070 1.405 ;
        END
        AntennaGateArea 0.0604 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.250 1.280 ;
        RECT  0.070 1.020 0.210 1.630 ;
        END
        AntennaGateArea 0.0413 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.020 0.790 1.375 ;
        END
        AntennaGateArea 0.0414 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.905 -0.210 1.680 0.210 ;
        RECT  0.735 -0.210 0.905 0.660 ;
        RECT  0.000 -0.210 0.735 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.585 2.310 1.680 2.730 ;
        RECT  1.415 1.775 1.585 2.730 ;
        RECT  0.805 2.310 1.415 2.730 ;
        RECT  0.115 2.015 0.805 2.730 ;
        RECT  0.000 2.310 0.115 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.310 1.050 1.370 1.310 ;
        RECT  1.190 0.780 1.310 1.310 ;
        RECT  0.490 0.780 1.190 0.900 ;
        RECT  0.490 1.585 0.555 1.755 ;
        RECT  0.370 0.780 0.490 1.755 ;
        RECT  0.265 0.780 0.370 0.900 ;
        RECT  0.095 0.730 0.265 0.900 ;
    END
END OAI2BB1XLAD
MACRO OAI2BB2X1AD
    CLASS CORE ;
    FOREIGN OAI2BB2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.600 2.170 1.725 ;
        RECT  2.000 0.600 2.030 0.860 ;
        RECT  1.725 1.605 2.030 1.725 ;
        RECT  1.555 1.605 1.725 2.035 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 1.105 1.330 1.395 ;
        END
        AntennaGateArea 0.09 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.105 1.625 1.485 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.140 0.925 1.375 ;
        END
        AntennaGateArea 0.041 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.000 0.270 1.260 ;
        RECT  0.070 0.585 0.210 1.260 ;
        END
        AntennaGateArea 0.0414 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.520 -0.210 2.240 0.210 ;
        RECT  1.260 -0.210 1.520 0.745 ;
        RECT  0.255 -0.210 1.260 0.210 ;
        RECT  0.085 -0.210 0.255 0.420 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.085 2.310 2.240 2.730 ;
        RECT  1.915 1.855 2.085 2.730 ;
        RECT  1.115 2.310 1.915 2.730 ;
        RECT  0.945 1.610 1.115 2.730 ;
        RECT  0.265 2.310 0.945 2.730 ;
        RECT  0.095 1.900 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.880 1.000 1.910 1.260 ;
        RECT  1.760 0.865 1.880 1.260 ;
        RECT  0.835 0.865 1.760 0.985 ;
        RECT  0.665 0.685 0.835 0.985 ;
        RECT  0.510 0.865 0.665 0.985 ;
        RECT  0.510 1.495 0.630 1.615 ;
        RECT  0.390 0.865 0.510 1.615 ;
        RECT  0.360 1.495 0.390 1.615 ;
    END
END OAI2BB2X1AD
MACRO OAI2BB2X2AD
    CLASS CORE ;
    FOREIGN OAI2BB2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 0.710 2.170 1.855 ;
        RECT  2.030 0.380 2.130 1.855 ;
        RECT  1.995 0.380 2.030 0.900 ;
        RECT  1.725 1.735 2.030 1.855 ;
        RECT  1.555 1.735 1.725 2.165 ;
        END
        AntennaDiffArea 0.401 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 1.020 1.330 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.020 1.625 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.120 0.925 1.375 ;
        END
        AntennaGateArea 0.075 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.000 0.270 1.260 ;
        RECT  0.070 0.585 0.210 1.260 ;
        END
        AntennaGateArea 0.0754 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.480 -0.210 2.240 0.210 ;
        RECT  1.220 -0.210 1.480 0.650 ;
        RECT  0.255 -0.210 1.220 0.210 ;
        RECT  0.085 -0.210 0.255 0.305 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.085 2.310 2.240 2.730 ;
        RECT  1.915 2.045 2.085 2.730 ;
        RECT  1.065 2.310 1.915 2.730 ;
        RECT  0.895 1.815 1.065 2.730 ;
        RECT  0.265 2.310 0.895 2.730 ;
        RECT  0.095 1.980 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.880 1.020 1.910 1.280 ;
        RECT  1.760 1.020 1.880 1.615 ;
        RECT  1.625 0.390 1.795 0.890 ;
        RECT  0.510 1.495 1.760 1.615 ;
        RECT  1.075 0.770 1.625 0.890 ;
        RECT  0.955 0.385 1.075 0.890 ;
        RECT  0.905 0.385 0.955 0.555 ;
        RECT  0.635 0.735 0.805 0.905 ;
        RECT  0.510 0.785 0.635 0.905 ;
        RECT  0.390 0.785 0.510 1.615 ;
        RECT  0.350 1.495 0.390 1.615 ;
    END
END OAI2BB2X2AD
MACRO OAI2BB2X4AD
    CLASS CORE ;
    FOREIGN OAI2BB2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.165 1.005 3.290 1.515 ;
        RECT  3.035 0.620 3.165 1.515 ;
        RECT  2.925 0.620 3.035 0.790 ;
        RECT  2.865 1.385 3.035 1.940 ;
        RECT  2.015 1.690 2.865 1.820 ;
        RECT  1.845 1.690 2.015 2.165 ;
        END
        AntennaDiffArea 0.664 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.110 2.580 1.230 ;
        RECT  2.320 1.110 2.440 1.570 ;
        RECT  1.535 1.450 2.320 1.570 ;
        RECT  1.415 1.110 1.535 1.570 ;
        RECT  1.190 1.110 1.415 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.110 2.200 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.705 1.110 1.050 1.375 ;
        END
        AntennaGateArea 0.144 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.225 0.985 0.345 1.375 ;
        RECT  0.070 1.145 0.225 1.375 ;
        END
        AntennaGateArea 0.144 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.375 -0.210 3.640 0.210 ;
        RECT  2.205 -0.210 2.375 0.510 ;
        RECT  1.625 -0.210 2.205 0.210 ;
        RECT  1.455 -0.210 1.625 0.485 ;
        RECT  0.275 -0.210 1.455 0.210 ;
        RECT  0.105 -0.210 0.275 0.785 ;
        RECT  0.000 -0.210 0.105 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.395 2.310 3.640 2.730 ;
        RECT  3.225 1.725 3.395 2.730 ;
        RECT  2.675 2.310 3.225 2.730 ;
        RECT  2.505 1.940 2.675 2.730 ;
        RECT  1.255 2.310 2.505 2.730 ;
        RECT  0.825 1.665 1.255 2.730 ;
        RECT  0.275 2.310 0.825 2.730 ;
        RECT  0.105 1.525 0.275 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  3.285 0.380 3.455 0.810 ;
        RECT  2.780 0.380 3.285 0.500 ;
        RECT  2.820 1.065 2.915 1.260 ;
        RECT  2.700 0.870 2.820 1.260 ;
        RECT  2.520 0.350 2.780 0.750 ;
        RECT  0.885 0.870 2.700 0.990 ;
        RECT  2.060 0.630 2.520 0.750 ;
        RECT  1.800 0.370 2.060 0.750 ;
        RECT  1.295 0.630 1.800 0.750 ;
        RECT  1.035 0.370 1.295 0.750 ;
        RECT  0.715 0.450 0.885 0.990 ;
        RECT  0.585 0.870 0.715 0.990 ;
        RECT  0.585 1.520 0.635 1.950 ;
        RECT  0.465 0.870 0.585 1.950 ;
    END
END OAI2BB2X4AD
MACRO OAI2BB2XLAD
    CLASS CORE ;
    FOREIGN OAI2BB2XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.555 2.170 1.725 ;
        RECT  2.000 0.555 2.030 0.815 ;
        RECT  1.725 1.605 2.030 1.725 ;
        RECT  1.555 1.605 1.725 1.775 ;
        END
        AntennaDiffArea 0.15 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 1.105 1.330 1.395 ;
        END
        AntennaGateArea 0.0604 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.105 1.625 1.485 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.140 0.925 1.375 ;
        END
        AntennaGateArea 0.041 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.000 0.270 1.260 ;
        RECT  0.070 0.585 0.210 1.260 ;
        END
        AntennaGateArea 0.0414 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.520 -0.210 2.240 0.210 ;
        RECT  1.260 -0.210 1.520 0.745 ;
        RECT  0.255 -0.210 1.260 0.210 ;
        RECT  0.085 -0.210 0.255 0.420 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.105 2.310 2.240 2.730 ;
        RECT  1.935 1.845 2.105 2.730 ;
        RECT  1.085 2.310 1.935 2.730 ;
        RECT  0.915 1.610 1.085 2.730 ;
        RECT  0.265 2.310 0.915 2.730 ;
        RECT  0.095 1.900 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.880 1.000 1.910 1.260 ;
        RECT  1.760 0.865 1.880 1.260 ;
        RECT  0.835 0.865 1.760 0.985 ;
        RECT  0.665 0.685 0.835 0.985 ;
        RECT  0.510 0.865 0.665 0.985 ;
        RECT  0.510 1.495 0.630 1.615 ;
        RECT  0.390 0.865 0.510 1.615 ;
        RECT  0.360 1.495 0.390 1.615 ;
    END
END OAI2BB2XLAD
MACRO OAI31X1AD
    CLASS CORE ;
    FOREIGN OAI31X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.690 1.610 1.655 ;
        RECT  1.425 0.690 1.470 0.860 ;
        RECT  1.175 1.525 1.470 1.655 ;
        RECT  1.005 1.525 1.175 1.955 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.020 1.350 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.230 1.265 ;
        END
        AntennaGateArea 0.09 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.005 0.700 1.265 ;
        RECT  0.490 1.145 0.580 1.265 ;
        RECT  0.350 1.145 0.490 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.020 1.050 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.855 -0.210 1.680 0.210 ;
        RECT  0.165 -0.210 0.855 0.385 ;
        RECT  0.000 -0.210 0.165 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.535 2.310 1.680 2.730 ;
        RECT  1.365 1.775 1.535 2.730 ;
        RECT  0.230 2.310 1.365 2.730 ;
        RECT  0.080 1.470 0.230 2.730 ;
        RECT  0.000 2.310 0.080 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.065 0.675 1.235 0.845 ;
        RECT  0.545 0.725 1.065 0.845 ;
        RECT  0.375 0.675 0.545 0.845 ;
    END
END OAI31X1AD
MACRO OAI31X2AD
    CLASS CORE ;
    FOREIGN OAI31X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.780 1.890 1.655 ;
        RECT  1.745 0.470 1.760 1.655 ;
        RECT  1.590 0.470 1.745 0.900 ;
        RECT  1.330 1.520 1.745 1.655 ;
        RECT  1.160 1.520 1.330 1.995 ;
        END
        AntennaDiffArea 0.401 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.040 1.625 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.235 1.050 0.505 1.265 ;
        RECT  0.130 1.050 0.235 1.375 ;
        RECT  0.070 1.145 0.130 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.055 0.900 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.020 1.050 1.330 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.040 -0.210 1.960 0.210 ;
        RECT  0.870 -0.210 1.040 0.675 ;
        RECT  0.320 -0.210 0.870 0.210 ;
        RECT  0.150 -0.210 0.320 0.840 ;
        RECT  0.000 -0.210 0.150 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.690 2.310 1.960 2.730 ;
        RECT  1.520 1.775 1.690 2.730 ;
        RECT  0.370 2.310 1.520 2.730 ;
        RECT  0.200 1.555 0.370 2.730 ;
        RECT  0.000 2.310 0.200 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.230 0.475 1.400 0.920 ;
        RECT  0.680 0.800 1.230 0.920 ;
        RECT  0.510 0.460 0.680 0.920 ;
    END
END OAI31X2AD
MACRO OAI31X4AD
    CLASS CORE ;
    FOREIGN OAI31X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.765 1.005 3.010 1.625 ;
        RECT  2.675 0.680 2.765 1.625 ;
        RECT  2.635 0.680 2.675 1.990 ;
        RECT  2.505 1.495 2.635 1.990 ;
        RECT  1.970 1.495 2.505 1.625 ;
        RECT  1.840 1.495 1.970 1.820 ;
        RECT  1.335 1.690 1.840 1.820 ;
        RECT  1.165 1.690 1.335 2.120 ;
        END
        AntennaDiffArea 0.664 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.015 2.500 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.015 0.860 2.135 1.275 ;
        RECT  0.510 0.860 2.015 0.980 ;
        RECT  0.390 0.860 0.510 1.375 ;
        RECT  0.325 1.050 0.390 1.375 ;
        RECT  0.070 1.145 0.325 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.110 1.860 1.230 ;
        RECT  1.600 1.110 1.720 1.570 ;
        RECT  0.900 1.450 1.600 1.570 ;
        RECT  0.630 1.100 0.900 1.570 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.090 1.100 1.480 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.055 -0.210 3.360 0.210 ;
        RECT  1.885 -0.210 2.055 0.500 ;
        RECT  1.335 -0.210 1.885 0.210 ;
        RECT  1.165 -0.210 1.335 0.500 ;
        RECT  0.615 -0.210 1.165 0.210 ;
        RECT  0.445 -0.210 0.615 0.500 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.035 2.310 3.360 2.730 ;
        RECT  2.865 1.845 3.035 2.730 ;
        RECT  2.315 2.310 2.865 2.730 ;
        RECT  2.145 1.800 2.315 2.730 ;
        RECT  0.375 2.310 2.145 2.730 ;
        RECT  0.205 1.515 0.375 2.730 ;
        RECT  0.000 2.310 0.205 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.970 0.440 3.140 0.870 ;
        RECT  2.465 0.440 2.970 0.560 ;
        RECT  2.205 0.360 2.465 0.740 ;
        RECT  1.740 0.620 2.205 0.740 ;
        RECT  1.480 0.360 1.740 0.740 ;
        RECT  1.020 0.620 1.480 0.740 ;
        RECT  0.760 0.360 1.020 0.740 ;
        RECT  0.255 0.620 0.760 0.740 ;
        RECT  0.085 0.365 0.255 0.795 ;
    END
END OAI31X4AD
MACRO OAI31XLAD
    CLASS CORE ;
    FOREIGN OAI31XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.735 1.610 1.655 ;
        RECT  1.425 0.735 1.470 0.905 ;
        RECT  1.175 1.525 1.470 1.655 ;
        RECT  1.005 1.525 1.175 1.720 ;
        END
        AntennaDiffArea 0.15 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.040 1.350 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.230 1.265 ;
        END
        AntennaGateArea 0.06 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 1.025 0.680 1.285 ;
        RECT  0.490 1.145 0.560 1.285 ;
        RECT  0.350 1.145 0.490 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 1.040 1.050 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.855 -0.210 1.680 0.210 ;
        RECT  0.165 -0.210 0.855 0.475 ;
        RECT  0.000 -0.210 0.165 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.580 2.310 1.680 2.730 ;
        RECT  1.320 1.775 1.580 2.730 ;
        RECT  0.255 2.310 1.320 2.730 ;
        RECT  0.085 1.645 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.065 0.735 1.235 0.905 ;
        RECT  0.545 0.785 1.065 0.905 ;
        RECT  0.375 0.735 0.545 0.905 ;
    END
END OAI31XLAD
MACRO OAI32X1AD
    CLASS CORE ;
    FOREIGN OAI32X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 1.030 1.890 1.630 ;
        RECT  1.730 0.650 1.850 1.630 ;
        RECT  1.575 0.650 1.730 0.820 ;
        RECT  1.335 1.510 1.730 1.630 ;
        RECT  1.165 1.510 1.335 1.940 ;
        END
        AntennaDiffArea 0.234 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.020 2.170 1.450 ;
        END
        AntennaGateArea 0.09 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.020 1.610 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.450 1.280 ;
        RECT  0.070 1.020 0.210 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 1.020 0.790 1.395 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.020 1.250 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.005 -0.210 2.240 0.210 ;
        RECT  0.835 -0.210 1.005 0.635 ;
        RECT  0.270 -0.210 0.835 0.210 ;
        RECT  0.110 -0.210 0.270 0.865 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.995 2.310 2.240 2.730 ;
        RECT  1.825 1.785 1.995 2.730 ;
        RECT  0.365 2.310 1.825 2.730 ;
        RECT  0.195 1.525 0.365 2.730 ;
        RECT  0.000 2.310 0.195 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.970 0.405 2.090 0.865 ;
        RECT  1.430 0.405 1.970 0.525 ;
        RECT  1.310 0.405 1.430 0.875 ;
        RECT  0.410 0.755 1.310 0.875 ;
    END
END OAI32X1AD
MACRO OAI32X2AD
    CLASS CORE ;
    FOREIGN OAI32X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 1.030 1.890 1.630 ;
        RECT  1.730 0.650 1.850 1.630 ;
        RECT  1.575 0.650 1.730 0.820 ;
        RECT  1.335 1.510 1.730 1.630 ;
        RECT  1.165 1.510 1.335 1.940 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.045 2.170 1.450 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.020 1.610 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.450 1.280 ;
        RECT  0.070 1.020 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.570 1.020 0.790 1.395 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.020 1.250 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.050 -0.210 2.240 0.210 ;
        RECT  0.790 -0.210 1.050 0.650 ;
        RECT  0.265 -0.210 0.790 0.210 ;
        RECT  0.095 -0.210 0.265 0.850 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.995 2.310 2.240 2.730 ;
        RECT  1.825 1.800 1.995 2.730 ;
        RECT  0.365 2.310 1.825 2.730 ;
        RECT  0.195 1.525 0.365 2.730 ;
        RECT  0.000 2.310 0.195 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.970 0.405 2.090 0.925 ;
        RECT  1.385 0.405 1.970 0.525 ;
        RECT  1.215 0.405 1.385 0.890 ;
        RECT  0.625 0.770 1.215 0.890 ;
        RECT  0.455 0.420 0.625 0.890 ;
    END
END OAI32X2AD
MACRO OAI32X4AD
    CLASS CORE ;
    FOREIGN OAI32X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.985 0.830 4.130 1.575 ;
        RECT  3.815 0.830 3.985 0.950 ;
        RECT  3.260 1.455 3.985 1.575 ;
        RECT  3.695 0.625 3.815 0.950 ;
        RECT  2.685 0.625 3.695 0.745 ;
        RECT  3.090 1.455 3.260 1.975 ;
        RECT  2.130 1.455 3.090 1.575 ;
        RECT  2.000 1.455 2.130 1.820 ;
        RECT  1.455 1.690 2.000 1.820 ;
        RECT  1.285 1.690 1.455 2.120 ;
        END
        AntennaDiffArea 0.89 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.575 1.090 3.825 1.210 ;
        RECT  3.455 0.865 3.575 1.210 ;
        RECT  2.730 0.865 3.455 0.985 ;
        RECT  2.590 0.865 2.730 1.260 ;
        END
        AntennaGateArea 0.324 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 1.110 3.335 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.150 0.860 2.270 1.275 ;
        RECT  0.510 0.860 2.150 0.980 ;
        RECT  0.390 0.860 0.510 1.375 ;
        RECT  0.340 1.005 0.390 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.110 2.010 1.230 ;
        RECT  1.750 1.110 1.870 1.570 ;
        RECT  0.770 1.450 1.750 1.570 ;
        RECT  0.770 1.110 0.990 1.230 ;
        RECT  0.630 1.110 0.770 1.570 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.375 1.100 1.630 1.220 ;
        RECT  1.110 1.100 1.375 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.175 -0.210 4.200 0.210 ;
        RECT  2.005 -0.210 2.175 0.500 ;
        RECT  1.455 -0.210 2.005 0.210 ;
        RECT  1.285 -0.210 1.455 0.500 ;
        RECT  0.735 -0.210 1.285 0.210 ;
        RECT  0.565 -0.210 0.735 0.500 ;
        RECT  0.000 -0.210 0.565 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.930 2.310 4.200 2.730 ;
        RECT  3.760 1.735 3.930 2.730 ;
        RECT  2.540 2.310 3.760 2.730 ;
        RECT  2.370 1.735 2.540 2.730 ;
        RECT  0.485 2.310 2.370 2.730 ;
        RECT  0.315 1.715 0.485 2.730 ;
        RECT  0.000 2.310 0.315 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  3.935 0.380 4.055 0.710 ;
        RECT  2.540 0.380 3.935 0.500 ;
        RECT  2.420 0.380 2.540 0.740 ;
        RECT  2.370 0.570 2.420 0.740 ;
        RECT  1.860 0.620 2.370 0.740 ;
        RECT  1.600 0.360 1.860 0.740 ;
        RECT  1.140 0.620 1.600 0.740 ;
        RECT  0.880 0.360 1.140 0.740 ;
        RECT  0.270 0.620 0.880 0.740 ;
        RECT  0.150 0.385 0.270 0.905 ;
    END
END OAI32X4AD
MACRO OAI32XLAD
    CLASS CORE ;
    FOREIGN OAI32XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.770 0.585 1.890 1.630 ;
        RECT  1.750 0.585 1.770 0.905 ;
        RECT  1.000 1.510 1.770 1.630 ;
        RECT  1.405 0.735 1.750 0.905 ;
        END
        AntennaDiffArea 0.156 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.025 1.650 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.020 1.350 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.370 1.280 ;
        RECT  0.070 1.020 0.210 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.560 1.020 0.770 1.380 ;
        END
        AntennaGateArea 0.06 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.885 1.110 2.005 ;
        RECT  0.350 1.705 0.490 2.005 ;
        END
        AntennaGateArea 0.06 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.795 -0.210 1.960 0.210 ;
        RECT  0.105 -0.210 0.795 0.475 ;
        RECT  0.000 -0.210 0.105 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.845 2.310 1.960 2.730 ;
        RECT  1.675 1.750 1.845 2.730 ;
        RECT  0.230 2.310 1.675 2.730 ;
        RECT  0.110 1.500 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.960 2.520 ;
        LAYER M1 ;
        RECT  1.260 0.330 1.565 0.450 ;
        RECT  1.045 0.330 1.260 0.880 ;
        RECT  0.330 0.760 1.045 0.880 ;
    END
END OAI32XLAD
MACRO OAI33X1AD
    CLASS CORE ;
    FOREIGN OAI33X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.595 2.450 1.655 ;
        RECT  2.185 0.385 2.310 0.765 ;
        RECT  1.275 1.525 2.310 1.655 ;
        RECT  1.680 0.385 2.185 0.505 ;
        RECT  1.560 0.385 1.680 0.680 ;
        RECT  1.420 0.560 1.560 0.680 ;
        RECT  1.105 1.525 1.275 1.955 ;
        END
        AntennaDiffArea 0.309 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.070 0.425 1.240 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.0906 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.705 0.770 1.935 ;
        RECT  0.585 1.040 0.730 1.935 ;
        END
        AntennaGateArea 0.09 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 1.040 1.070 1.375 ;
        END
        AntennaGateArea 0.0906 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.040 2.190 1.375 ;
        END
        AntennaGateArea 0.0906 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.615 1.040 1.890 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.070 1.475 1.375 ;
        END
        AntennaGateArea 0.09 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.815 -0.210 2.520 0.210 ;
        RECT  0.125 -0.210 0.815 0.385 ;
        RECT  0.000 -0.210 0.125 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.265 2.310 2.520 2.730 ;
        RECT  2.095 1.785 2.265 2.730 ;
        RECT  0.310 2.310 2.095 2.730 ;
        RECT  0.125 1.525 0.310 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.825 0.625 1.995 0.920 ;
        RECT  1.275 0.800 1.825 0.920 ;
        RECT  1.105 0.570 1.275 0.920 ;
        RECT  0.575 0.800 1.105 0.920 ;
        RECT  0.405 0.665 0.575 0.920 ;
    END
END OAI33X1AD
MACRO OAI33X2AD
    CLASS CORE ;
    FOREIGN OAI33X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.690 2.450 1.655 ;
        RECT  2.310 0.385 2.415 1.655 ;
        RECT  2.245 0.385 2.310 0.835 ;
        RECT  1.335 1.525 2.310 1.655 ;
        RECT  1.695 0.385 2.245 0.505 ;
        RECT  1.525 0.385 1.695 0.555 ;
        RECT  1.165 1.525 1.335 1.955 ;
        END
        AntennaDiffArea 0.581 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.065 0.425 1.235 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.775 1.705 0.815 1.935 ;
        RECT  0.630 1.020 0.775 1.935 ;
        END
        AntennaGateArea 0.162 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.895 1.020 1.070 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.020 2.190 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.615 1.020 1.890 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.020 1.475 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.020 -0.210 2.520 0.210 ;
        RECT  0.760 -0.210 1.020 0.650 ;
        RECT  0.255 -0.210 0.760 0.210 ;
        RECT  0.085 -0.210 0.255 0.730 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.295 2.310 2.520 2.730 ;
        RECT  2.125 1.845 2.295 2.730 ;
        RECT  0.350 2.310 2.125 2.730 ;
        RECT  0.165 1.525 0.350 2.730 ;
        RECT  0.000 2.310 0.165 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.885 0.625 2.055 0.900 ;
        RECT  1.335 0.780 1.885 0.900 ;
        RECT  1.165 0.405 1.335 0.900 ;
        RECT  0.615 0.780 1.165 0.900 ;
        RECT  0.445 0.405 0.615 0.900 ;
    END
END OAI33X2AD
MACRO OAI33X4AD
    CLASS CORE ;
    FOREIGN OAI33X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 0.770 4.690 1.820 ;
        RECT  4.360 0.770 4.550 0.900 ;
        RECT  3.595 1.690 4.550 1.820 ;
        RECT  4.240 0.625 4.360 0.900 ;
        RECT  2.660 0.625 4.240 0.745 ;
        RECT  3.425 1.690 3.595 2.135 ;
        RECT  1.435 1.690 3.425 1.820 ;
        RECT  1.265 1.690 1.435 2.120 ;
        END
        AntennaDiffArea 1.024 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.105 0.860 2.225 1.275 ;
        RECT  0.510 0.860 2.105 0.980 ;
        RECT  0.390 0.860 0.510 1.375 ;
        RECT  0.350 1.025 0.390 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.845 1.120 1.960 1.240 ;
        RECT  1.725 1.120 1.845 1.570 ;
        RECT  1.700 1.120 1.725 1.240 ;
        RECT  1.000 1.450 1.725 1.570 ;
        RECT  0.880 1.100 1.000 1.570 ;
        RECT  0.630 1.100 0.880 1.380 ;
        END
        AntennaGateArea 0.324 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.145 1.100 1.460 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.260 1.020 4.380 1.570 ;
        RECT  2.750 1.450 4.260 1.570 ;
        RECT  2.590 1.015 2.750 1.570 ;
        END
        AntennaGateArea 0.324 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.960 0.865 4.080 1.280 ;
        RECT  3.110 0.865 3.960 0.985 ;
        RECT  2.870 0.865 3.110 1.260 ;
        END
        AntennaGateArea 0.324 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 1.110 3.760 1.330 ;
        END
        AntennaGateArea 0.324 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.155 -0.210 4.760 0.210 ;
        RECT  1.985 -0.210 2.155 0.485 ;
        RECT  1.435 -0.210 1.985 0.210 ;
        RECT  1.265 -0.210 1.435 0.485 ;
        RECT  0.715 -0.210 1.265 0.210 ;
        RECT  0.545 -0.210 0.715 0.485 ;
        RECT  0.000 -0.210 0.545 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.555 2.310 4.760 2.730 ;
        RECT  4.385 1.990 4.555 2.730 ;
        RECT  2.585 2.310 4.385 2.730 ;
        RECT  2.415 1.975 2.585 2.730 ;
        RECT  0.475 2.310 2.415 2.730 ;
        RECT  0.305 1.555 0.475 2.730 ;
        RECT  0.000 2.310 0.305 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.760 2.520 ;
        LAYER M1 ;
        RECT  4.505 0.380 4.675 0.550 ;
        RECT  2.515 0.380 4.505 0.500 ;
        RECT  2.345 0.355 2.515 0.785 ;
        RECT  1.795 0.620 2.345 0.740 ;
        RECT  1.625 0.505 1.795 0.740 ;
        RECT  1.075 0.620 1.625 0.740 ;
        RECT  0.905 0.500 1.075 0.740 ;
        RECT  0.400 0.620 0.905 0.740 ;
        RECT  0.140 0.360 0.400 0.740 ;
    END
END OAI33X4AD
MACRO OAI33XLAD
    CLASS CORE ;
    FOREIGN OAI33XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.735 2.450 1.655 ;
        RECT  2.310 0.520 2.350 1.655 ;
        RECT  2.225 0.520 2.310 0.905 ;
        RECT  1.275 1.525 2.310 1.655 ;
        RECT  1.440 0.520 2.225 0.640 ;
        RECT  1.105 1.525 1.275 1.695 ;
        END
        AntennaDiffArea 0.264 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.065 0.425 1.235 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.705 0.770 1.935 ;
        RECT  0.585 1.020 0.730 1.935 ;
        END
        AntennaGateArea 0.06 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 1.020 1.070 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.020 2.190 1.375 ;
        END
        AntennaGateArea 0.0604 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.615 1.020 1.890 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.070 1.475 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.815 -0.210 2.520 0.210 ;
        RECT  0.125 -0.210 0.815 0.475 ;
        RECT  0.000 -0.210 0.125 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.295 2.310 2.520 2.730 ;
        RECT  2.125 1.775 2.295 2.730 ;
        RECT  0.310 2.310 2.125 2.730 ;
        RECT  0.125 1.525 0.310 2.730 ;
        RECT  0.000 2.310 0.125 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  0.360 0.760 2.080 0.880 ;
    END
END OAI33XLAD
MACRO OR2X1AD
    CLASS CORE ;
    FOREIGN OR2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.305 0.650 1.330 1.375 ;
        RECT  1.160 0.650 1.305 1.835 ;
        RECT  1.135 1.405 1.160 1.835 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.015 0.770 1.375 ;
        END
        AntennaGateArea 0.0563 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.240 1.260 ;
        END
        AntennaGateArea 0.056 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.925 -0.210 1.400 0.210 ;
        RECT  0.755 -0.210 0.925 0.475 ;
        RECT  0.255 -0.210 0.755 0.210 ;
        RECT  0.085 -0.210 0.255 0.470 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 2.310 1.400 2.730 ;
        RECT  0.775 1.525 0.945 2.730 ;
        RECT  0.000 2.310 0.775 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.920 0.760 1.040 1.280 ;
        RECT  0.480 0.760 0.920 0.880 ;
        RECT  0.360 0.760 0.480 1.600 ;
        RECT  0.095 1.430 0.360 1.600 ;
    END
END OR2X1AD
MACRO OR2X2AD
    CLASS CORE ;
    FOREIGN OR2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 0.865 1.330 1.375 ;
        RECT  1.170 0.420 1.290 2.020 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 0.980 0.770 1.375 ;
        END
        AntennaGateArea 0.0924 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.230 1.260 ;
        END
        AntennaGateArea 0.092 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.885 -0.210 1.400 0.210 ;
        RECT  0.715 -0.210 0.885 0.375 ;
        RECT  0.270 -0.210 0.715 0.210 ;
        RECT  0.100 -0.210 0.270 0.375 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.955 2.310 1.400 2.730 ;
        RECT  0.785 1.545 0.955 2.730 ;
        RECT  0.000 2.310 0.785 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.930 0.725 1.050 1.280 ;
        RECT  0.475 0.725 0.930 0.845 ;
        RECT  0.355 0.725 0.475 1.625 ;
        RECT  0.275 1.455 0.355 1.625 ;
        RECT  0.105 1.455 0.275 1.885 ;
    END
END OR2X2AD
MACRO OR2X4AD
    CLASS CORE ;
    FOREIGN OR2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.730 2.170 1.515 ;
        RECT  1.965 0.730 2.030 0.860 ;
        RECT  1.965 1.385 2.030 1.515 ;
        RECT  1.795 0.415 1.965 0.860 ;
        RECT  1.795 1.385 1.965 2.130 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.265 1.035 1.385 1.570 ;
        RECT  0.490 1.450 1.265 1.570 ;
        RECT  0.255 1.160 0.490 1.655 ;
        END
        AntennaGateArea 0.1842 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.615 1.080 1.135 1.330 ;
        END
        AntennaGateArea 0.184 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.325 -0.210 2.520 0.210 ;
        RECT  2.155 -0.210 2.325 0.565 ;
        RECT  1.605 -0.210 2.155 0.210 ;
        RECT  1.435 -0.210 1.605 0.565 ;
        RECT  0.885 -0.210 1.435 0.210 ;
        RECT  0.715 -0.210 0.885 0.825 ;
        RECT  0.000 -0.210 0.715 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.325 2.310 2.520 2.730 ;
        RECT  2.155 1.690 2.325 2.730 ;
        RECT  1.605 2.310 2.155 2.730 ;
        RECT  1.435 1.995 1.605 2.730 ;
        RECT  0.310 2.310 1.435 2.730 ;
        RECT  0.140 1.795 0.310 2.730 ;
        RECT  0.000 2.310 0.140 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  1.665 1.075 1.890 1.245 ;
        RECT  1.545 0.725 1.665 1.875 ;
        RECT  1.245 0.725 1.545 0.845 ;
        RECT  0.940 1.730 1.545 1.875 ;
        RECT  1.075 0.395 1.245 0.845 ;
        RECT  0.770 1.730 0.940 2.160 ;
    END
END OR2X4AD
MACRO OR2X6AD
    CLASS CORE ;
    FOREIGN OR2X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 0.395 2.715 0.825 ;
        RECT  2.545 1.415 2.715 2.145 ;
        RECT  2.510 0.645 2.545 0.825 ;
        RECT  2.510 1.415 2.545 1.655 ;
        RECT  2.310 0.645 2.510 1.655 ;
        RECT  1.995 0.645 2.310 0.825 ;
        RECT  1.995 1.415 2.310 1.655 ;
        RECT  1.825 0.385 1.995 0.825 ;
        RECT  1.825 1.415 1.995 2.145 ;
        END
        AntennaDiffArea 0.795 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.335 1.080 1.405 1.250 ;
        RECT  1.215 1.080 1.335 1.570 ;
        RECT  0.640 1.450 1.215 1.570 ;
        RECT  0.500 1.085 0.640 1.570 ;
        RECT  0.255 1.085 0.500 1.380 ;
        RECT  0.240 1.085 0.255 1.255 ;
        END
        AntennaGateArea 0.2689 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 1.080 1.095 1.330 ;
        END
        AntennaGateArea 0.2673 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.355 -0.210 2.800 0.210 ;
        RECT  2.185 -0.210 2.355 0.510 ;
        RECT  1.635 -0.210 2.185 0.210 ;
        RECT  1.465 -0.210 1.635 0.575 ;
        RECT  0.865 -0.210 1.465 0.210 ;
        RECT  0.695 -0.210 0.865 0.465 ;
        RECT  0.275 -0.210 0.695 0.210 ;
        RECT  0.105 -0.210 0.275 0.465 ;
        RECT  0.000 -0.210 0.105 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.355 2.310 2.800 2.730 ;
        RECT  2.185 1.840 2.355 2.730 ;
        RECT  1.575 2.310 2.185 2.730 ;
        RECT  1.405 1.965 1.575 2.730 ;
        RECT  0.290 2.310 1.405 2.730 ;
        RECT  0.120 1.685 0.290 2.730 ;
        RECT  0.000 2.310 0.120 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  1.655 1.100 2.185 1.220 ;
        RECT  1.535 0.735 1.655 1.810 ;
        RECT  1.255 0.735 1.535 0.905 ;
        RECT  0.925 1.690 1.535 1.810 ;
        RECT  1.085 0.385 1.255 0.905 ;
        RECT  0.415 0.735 1.085 0.905 ;
        RECT  0.755 1.690 0.925 2.125 ;
    END
END OR2X6AD
MACRO OR2X8AD
    CLASS CORE ;
    FOREIGN OR2X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.005 0.415 3.175 2.155 ;
        RECT  2.730 0.630 3.005 1.700 ;
        RECT  2.455 0.630 2.730 0.895 ;
        RECT  2.455 1.365 2.730 1.700 ;
        RECT  2.285 0.385 2.455 0.895 ;
        RECT  2.285 1.365 2.455 2.155 ;
        END
        AntennaDiffArea 0.844 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 1.030 1.920 1.450 ;
        RECT  1.030 1.330 1.800 1.450 ;
        RECT  0.510 1.140 1.030 1.450 ;
        END
        AntennaGateArea 0.3707 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.035 1.680 1.210 ;
        RECT  1.160 0.900 1.280 1.210 ;
        RECT  0.390 0.900 1.160 1.020 ;
        RECT  0.270 0.900 0.390 1.375 ;
        RECT  0.070 1.145 0.270 1.375 ;
        END
        AntennaGateArea 0.369 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.535 -0.210 3.640 0.210 ;
        RECT  3.365 -0.210 3.535 0.830 ;
        RECT  2.815 -0.210 3.365 0.210 ;
        RECT  2.645 -0.210 2.815 0.490 ;
        RECT  2.095 -0.210 2.645 0.210 ;
        RECT  1.925 -0.210 2.095 0.645 ;
        RECT  1.360 -0.210 1.925 0.210 ;
        RECT  0.840 -0.210 1.360 0.540 ;
        RECT  0.265 -0.210 0.840 0.210 ;
        RECT  0.095 -0.210 0.265 0.720 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.535 2.310 3.640 2.730 ;
        RECT  3.365 1.465 3.535 2.730 ;
        RECT  2.815 2.310 3.365 2.730 ;
        RECT  2.645 1.845 2.815 2.730 ;
        RECT  2.095 2.310 2.645 2.730 ;
        RECT  1.925 1.845 2.095 2.730 ;
        RECT  0.875 2.310 1.925 2.730 ;
        RECT  0.705 1.845 0.875 2.730 ;
        RECT  0.000 2.310 0.705 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  2.160 1.050 2.600 1.220 ;
        RECT  2.040 0.785 2.160 1.690 ;
        RECT  1.735 0.785 2.040 0.905 ;
        RECT  1.485 1.570 2.040 1.690 ;
        RECT  1.565 0.475 1.735 0.905 ;
        RECT  0.625 0.660 1.565 0.780 ;
        RECT  1.315 1.570 1.485 2.000 ;
        RECT  0.265 1.570 1.315 1.690 ;
        RECT  0.455 0.550 0.625 0.780 ;
        RECT  0.095 1.570 0.265 2.000 ;
    END
END OR2X8AD
MACRO OR2XLAD
    CLASS CORE ;
    FOREIGN OR2XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 0.690 1.330 1.705 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.015 0.770 1.375 ;
        END
        AntennaGateArea 0.0444 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.240 1.260 ;
        END
        AntennaGateArea 0.044 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.925 -0.210 1.400 0.210 ;
        RECT  0.755 -0.210 0.925 0.475 ;
        RECT  0.255 -0.210 0.755 0.210 ;
        RECT  0.085 -0.210 0.255 0.470 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.945 2.310 1.400 2.730 ;
        RECT  0.775 1.575 0.945 2.730 ;
        RECT  0.000 2.310 0.775 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.400 2.520 ;
        LAYER M1 ;
        RECT  0.920 0.760 1.040 1.280 ;
        RECT  0.480 0.760 0.920 0.880 ;
        RECT  0.360 0.760 0.480 1.580 ;
        RECT  0.095 1.410 0.360 1.580 ;
    END
END OR2XLAD
MACRO OR3X1AD
    CLASS CORE ;
    FOREIGN OR3X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.640 1.610 1.920 ;
        RECT  1.410 0.640 1.470 0.900 ;
        RECT  1.440 1.400 1.470 1.920 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.015 1.050 1.490 ;
        END
        AntennaGateArea 0.073 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.000 0.775 1.660 ;
        END
        AntennaGateArea 0.073 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 1.025 0.270 1.285 ;
        RECT  0.110 1.025 0.240 1.375 ;
        RECT  0.070 1.145 0.110 1.375 ;
        END
        AntennaGateArea 0.0735 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.215 -0.210 1.680 0.210 ;
        RECT  1.045 -0.210 1.215 0.475 ;
        RECT  0.635 -0.210 1.045 0.210 ;
        RECT  0.465 -0.210 0.635 0.475 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.235 2.310 1.680 2.730 ;
        RECT  1.065 1.705 1.235 2.730 ;
        RECT  0.000 2.310 1.065 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.290 1.020 1.350 1.280 ;
        RECT  1.170 0.760 1.290 1.280 ;
        RECT  0.510 0.760 1.170 0.880 ;
        RECT  0.390 0.760 0.510 1.615 ;
        RECT  0.255 0.760 0.390 0.880 ;
        RECT  0.285 1.495 0.390 1.615 ;
        RECT  0.115 1.495 0.285 1.665 ;
        RECT  0.085 0.735 0.255 0.905 ;
    END
END OR3X1AD
MACRO OR3X2AD
    CLASS CORE ;
    FOREIGN OR3X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.350 1.610 2.075 ;
        RECT  1.440 0.350 1.470 0.870 ;
        RECT  1.440 1.555 1.470 2.075 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.015 1.060 1.465 ;
        END
        AntennaGateArea 0.12 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.000 0.770 1.660 ;
        END
        AntennaGateArea 0.12 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 1.025 0.270 1.285 ;
        RECT  0.110 1.025 0.240 1.375 ;
        RECT  0.070 1.145 0.110 1.375 ;
        END
        AntennaGateArea 0.12 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.165 -0.210 1.680 0.210 ;
        RECT  0.995 -0.210 1.165 0.390 ;
        RECT  0.635 -0.210 0.995 0.210 ;
        RECT  0.465 -0.210 0.635 0.390 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.235 2.310 1.680 2.730 ;
        RECT  1.065 1.600 1.235 2.730 ;
        RECT  0.000 2.310 1.065 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.305 1.020 1.350 1.280 ;
        RECT  1.185 0.725 1.305 1.280 ;
        RECT  0.510 0.725 1.185 0.845 ;
        RECT  0.390 0.725 0.510 1.720 ;
        RECT  0.255 0.725 0.390 0.845 ;
        RECT  0.285 1.600 0.390 1.720 ;
        RECT  0.115 1.600 0.285 2.030 ;
        RECT  0.085 0.700 0.255 0.870 ;
    END
END OR3X2AD
MACRO OR3X4AD
    CLASS CORE ;
    FOREIGN OR3X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 1.005 2.450 1.515 ;
        RECT  2.220 0.360 2.350 1.965 ;
        RECT  2.190 0.360 2.220 0.880 ;
        RECT  2.165 1.535 2.220 1.965 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.020 1.800 1.570 ;
        RECT  0.420 1.450 1.680 1.570 ;
        RECT  0.300 1.140 0.420 1.570 ;
        RECT  0.070 1.140 0.300 1.375 ;
        END
        AntennaGateArea 0.24 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 0.900 1.530 1.020 ;
        RECT  0.350 0.585 0.490 1.020 ;
        END
        AntennaGateArea 0.24 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.780 1.140 1.150 1.330 ;
        END
        AntennaGateArea 0.24 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.695 -0.210 2.800 0.210 ;
        RECT  2.525 -0.210 2.695 0.795 ;
        RECT  1.975 -0.210 2.525 0.210 ;
        RECT  1.805 -0.210 1.975 0.470 ;
        RECT  1.235 -0.210 1.805 0.210 ;
        RECT  1.065 -0.210 1.235 0.470 ;
        RECT  0.000 -0.210 1.065 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.695 2.310 2.800 2.730 ;
        RECT  2.525 1.715 2.695 2.730 ;
        RECT  1.975 2.310 2.525 2.730 ;
        RECT  1.805 1.995 1.975 2.730 ;
        RECT  0.255 2.310 1.805 2.730 ;
        RECT  0.085 1.730 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.040 1.020 2.100 1.280 ;
        RECT  1.920 0.620 2.040 1.830 ;
        RECT  1.660 0.620 1.920 0.740 ;
        RECT  1.115 1.710 1.920 1.830 ;
        RECT  1.400 0.340 1.660 0.740 ;
        RECT  0.910 0.620 1.400 0.740 ;
        RECT  0.945 1.710 1.115 2.140 ;
        RECT  0.650 0.340 0.910 0.740 ;
    END
END OR3X4AD
MACRO OR3X6AD
    CLASS CORE ;
    FOREIGN OR3X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.905 0.360 4.085 0.900 ;
        RECT  3.905 1.475 4.075 2.165 ;
        RECT  3.900 0.720 3.905 0.900 ;
        RECT  3.900 1.475 3.905 1.655 ;
        RECT  3.660 0.720 3.900 1.655 ;
        RECT  3.420 0.720 3.660 0.900 ;
        RECT  3.365 1.475 3.660 1.655 ;
        RECT  3.240 0.360 3.420 0.900 ;
        RECT  3.185 1.475 3.365 2.165 ;
        END
        AntennaDiffArea 0.795 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.700 1.040 2.820 1.570 ;
        RECT  1.330 1.450 2.700 1.570 ;
        RECT  1.190 1.110 1.330 1.570 ;
        RECT  1.060 1.110 1.190 1.230 ;
        END
        AntennaGateArea 0.361 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.370 0.870 2.490 1.260 ;
        RECT  1.590 0.870 2.370 0.990 ;
        RECT  1.470 0.870 1.590 1.280 ;
        RECT  0.680 0.870 1.470 0.990 ;
        RECT  0.560 0.870 0.680 1.330 ;
        RECT  0.305 1.190 0.560 1.330 ;
        END
        AntennaGateArea 0.361 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 1.140 2.215 1.330 ;
        END
        AntennaGateArea 0.361 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.745 -0.210 4.200 0.210 ;
        RECT  3.575 -0.210 3.745 0.580 ;
        RECT  3.000 -0.210 3.575 0.210 ;
        RECT  2.740 -0.210 3.000 0.240 ;
        RECT  2.265 -0.210 2.740 0.210 ;
        RECT  2.005 -0.210 2.265 0.510 ;
        RECT  1.325 -0.210 2.005 0.210 ;
        RECT  1.065 -0.210 1.325 0.510 ;
        RECT  0.255 -0.210 1.065 0.210 ;
        RECT  0.085 -0.210 0.255 0.765 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.715 2.310 4.200 2.730 ;
        RECT  3.545 1.845 3.715 2.730 ;
        RECT  2.995 2.310 3.545 2.730 ;
        RECT  2.825 1.935 2.995 2.730 ;
        RECT  1.155 2.310 2.825 2.730 ;
        RECT  0.985 1.935 1.155 2.730 ;
        RECT  0.000 2.310 0.985 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  3.065 1.065 3.505 1.235 ;
        RECT  2.945 0.630 3.065 1.810 ;
        RECT  0.480 0.630 2.945 0.750 ;
        RECT  2.065 1.690 2.945 1.810 ;
        RECT  1.895 1.690 2.065 2.120 ;
        RECT  0.255 1.690 1.895 1.810 ;
        RECT  0.085 1.690 0.255 2.120 ;
    END
END OR3X6AD
MACRO OR3X8AD
    CLASS CORE ;
    FOREIGN OR3X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.820 0.365 5.020 2.160 ;
        RECT  4.305 1.005 4.820 1.515 ;
        RECT  4.105 0.365 4.305 2.155 ;
        END
        AntennaDiffArea 0.844 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.560 1.020 3.680 1.620 ;
        RECT  2.170 1.500 3.560 1.620 ;
        RECT  1.910 1.140 2.170 1.620 ;
        RECT  0.490 1.500 1.910 1.620 ;
        RECT  0.375 1.145 0.490 1.620 ;
        RECT  0.350 1.065 0.375 1.620 ;
        RECT  0.205 1.065 0.350 1.285 ;
        END
        AntennaGateArea 0.48 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.260 1.020 3.380 1.380 ;
        RECT  2.470 1.260 3.260 1.380 ;
        RECT  2.350 0.900 2.470 1.380 ;
        RECT  1.610 0.900 2.350 1.020 ;
        RECT  1.490 0.900 1.610 1.380 ;
        RECT  1.405 0.980 1.490 1.380 ;
        RECT  0.730 1.260 1.405 1.380 ;
        RECT  0.610 0.790 0.730 1.380 ;
        RECT  0.570 0.790 0.610 1.050 ;
        END
        AntennaGateArea 0.48 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.020 2.990 1.140 ;
        RECT  2.730 0.660 2.850 1.140 ;
        RECT  1.250 0.660 2.730 0.780 ;
        RECT  1.130 0.660 1.250 1.140 ;
        RECT  0.910 0.865 1.130 1.140 ;
        END
        AntennaGateArea 0.48 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.365 -0.210 5.600 0.210 ;
        RECT  5.195 -0.210 5.365 0.795 ;
        RECT  4.645 -0.210 5.195 0.210 ;
        RECT  4.475 -0.210 4.645 0.795 ;
        RECT  3.915 -0.210 4.475 0.210 ;
        RECT  3.745 -0.210 3.915 0.645 ;
        RECT  3.115 -0.210 3.745 0.210 ;
        RECT  2.855 -0.210 3.115 0.250 ;
        RECT  1.920 -0.210 2.855 0.210 ;
        RECT  1.660 -0.210 1.920 0.250 ;
        RECT  1.005 -0.210 1.660 0.210 ;
        RECT  0.835 -0.210 1.005 0.645 ;
        RECT  0.000 -0.210 0.835 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.365 2.310 5.600 2.730 ;
        RECT  5.195 1.465 5.365 2.730 ;
        RECT  4.635 2.310 5.195 2.730 ;
        RECT  4.465 1.725 4.635 2.730 ;
        RECT  3.925 2.310 4.465 2.730 ;
        RECT  3.665 1.980 3.925 2.730 ;
        RECT  2.080 2.310 3.665 2.730 ;
        RECT  1.820 1.980 2.080 2.730 ;
        RECT  0.230 2.310 1.820 2.730 ;
        RECT  0.110 1.530 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  3.920 1.000 3.980 1.260 ;
        RECT  3.800 0.780 3.920 1.860 ;
        RECT  3.600 0.780 3.800 0.900 ;
        RECT  3.000 1.740 3.800 1.860 ;
        RECT  3.460 0.460 3.600 0.900 ;
        RECT  3.340 0.420 3.460 0.900 ;
        RECT  1.150 0.420 3.340 0.540 ;
        RECT  2.740 1.740 3.000 2.120 ;
        RECT  1.160 1.740 2.740 1.860 ;
        RECT  0.900 1.740 1.160 2.120 ;
    END
END OR3X8AD
MACRO OR3XLAD
    CLASS CORE ;
    FOREIGN OR3XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.735 1.610 1.665 ;
        RECT  1.425 0.735 1.470 0.905 ;
        RECT  1.425 1.495 1.470 1.665 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.015 1.060 1.415 ;
        END
        AntennaGateArea 0.056 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.000 0.770 1.660 ;
        END
        AntennaGateArea 0.056 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 1.025 0.270 1.285 ;
        RECT  0.110 1.025 0.240 1.375 ;
        RECT  0.070 1.145 0.110 1.375 ;
        END
        AntennaGateArea 0.0564 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.215 -0.210 1.680 0.210 ;
        RECT  1.045 -0.210 1.215 0.475 ;
        RECT  0.635 -0.210 1.045 0.210 ;
        RECT  0.465 -0.210 0.635 0.475 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.235 2.310 1.680 2.730 ;
        RECT  1.065 1.540 1.235 2.730 ;
        RECT  0.000 2.310 1.065 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 1.680 2.520 ;
        LAYER M1 ;
        RECT  1.305 1.020 1.350 1.280 ;
        RECT  1.185 0.760 1.305 1.280 ;
        RECT  0.510 0.760 1.185 0.880 ;
        RECT  0.390 0.760 0.510 1.615 ;
        RECT  0.255 0.760 0.390 0.880 ;
        RECT  0.285 1.495 0.390 1.615 ;
        RECT  0.115 1.495 0.285 1.665 ;
        RECT  0.085 0.735 0.255 0.905 ;
    END
END OR3XLAD
MACRO OR4X1AD
    CLASS CORE ;
    FOREIGN OR4X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.140 2.170 1.375 ;
        RECT  2.000 0.620 2.120 1.860 ;
        END
        AntennaDiffArea 0.207 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.000 1.640 1.440 ;
        END
        AntennaGateArea 0.065 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.020 1.330 1.375 ;
        END
        AntennaGateArea 0.065 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.000 0.820 1.465 ;
        END
        AntennaGateArea 0.065 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.000 0.490 1.465 ;
        END
        AntennaGateArea 0.0655 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.210 2.240 0.210 ;
        RECT  1.595 -0.210 1.765 0.640 ;
        RECT  0.995 -0.210 1.595 0.210 ;
        RECT  0.825 -0.210 0.995 0.470 ;
        RECT  0.255 -0.210 0.825 0.210 ;
        RECT  0.085 -0.210 0.255 0.640 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.750 2.310 2.240 2.730 ;
        RECT  1.580 1.575 1.750 2.730 ;
        RECT  0.000 2.310 1.580 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.760 0.760 1.880 1.280 ;
        RECT  0.230 0.760 1.760 0.880 ;
        RECT  0.230 1.600 0.365 1.770 ;
        RECT  0.110 0.760 0.230 1.770 ;
    END
END OR4X1AD
MACRO OR4X2AD
    CLASS CORE ;
    FOREIGN OR4X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.130 1.140 2.170 1.375 ;
        RECT  2.010 0.420 2.130 2.010 ;
        RECT  1.930 1.490 2.010 2.010 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.000 1.640 1.435 ;
        END
        AntennaGateArea 0.1103 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.020 1.330 1.375 ;
        END
        AntennaGateArea 0.11 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.000 0.820 1.465 ;
        END
        AntennaGateArea 0.11 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.020 0.510 1.465 ;
        END
        AntennaGateArea 0.11 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.795 -0.210 2.240 0.210 ;
        RECT  1.625 -0.210 1.795 0.605 ;
        RECT  1.025 -0.210 1.625 0.210 ;
        RECT  0.855 -0.210 1.025 0.640 ;
        RECT  0.255 -0.210 0.855 0.210 ;
        RECT  0.085 -0.210 0.255 0.640 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.685 2.310 2.240 2.730 ;
        RECT  1.515 1.595 1.685 2.730 ;
        RECT  0.000 2.310 1.515 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.760 0.760 1.880 1.280 ;
        RECT  0.230 0.760 1.760 0.880 ;
        RECT  0.230 1.595 0.395 2.025 ;
        RECT  0.110 0.760 0.230 2.025 ;
    END
END OR4X2AD
MACRO OR4X4AD
    CLASS CORE ;
    FOREIGN OR4X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.975 0.385 3.010 1.515 ;
        RECT  2.855 0.385 2.975 1.985 ;
        RECT  2.815 0.385 2.855 0.815 ;
        RECT  2.735 1.555 2.855 1.985 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.020 2.360 1.530 ;
        RECT  2.040 1.410 2.240 1.530 ;
        RECT  1.920 1.410 2.040 1.810 ;
        RECT  0.380 1.690 1.920 1.810 ;
        RECT  0.260 1.085 0.380 1.810 ;
        RECT  0.205 1.085 0.260 1.375 ;
        RECT  0.070 1.145 0.205 1.375 ;
        END
        AntennaGateArea 0.2188 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.940 1.020 2.060 1.290 ;
        RECT  1.800 1.170 1.940 1.290 ;
        RECT  1.680 1.170 1.800 1.570 ;
        RECT  0.770 1.450 1.680 1.570 ;
        RECT  0.630 1.145 0.770 1.570 ;
        RECT  0.510 0.710 0.630 1.570 ;
        END
        AntennaGateArea 0.218 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.095 0.900 1.780 1.020 ;
        RECT  0.820 0.630 1.095 1.020 ;
        END
        AntennaGateArea 0.218 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 1.190 1.420 1.330 ;
        RECT  1.030 1.140 1.290 1.330 ;
        RECT  0.975 1.190 1.030 1.330 ;
        END
        AntennaGateArea 0.218 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.345 -0.210 3.640 0.210 ;
        RECT  3.175 -0.210 3.345 0.815 ;
        RECT  2.670 -0.210 3.175 0.210 ;
        RECT  2.410 -0.210 2.670 0.575 ;
        RECT  1.920 -0.210 2.410 0.210 ;
        RECT  1.660 -0.210 1.920 0.540 ;
        RECT  1.200 -0.210 1.660 0.210 ;
        RECT  0.940 -0.210 1.200 0.500 ;
        RECT  0.000 -0.210 0.940 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.265 2.310 3.640 2.730 ;
        RECT  3.095 1.735 3.265 2.730 ;
        RECT  2.570 2.310 3.095 2.730 ;
        RECT  2.400 1.890 2.570 2.730 ;
        RECT  0.255 2.310 2.400 2.730 ;
        RECT  0.085 1.995 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  2.615 0.995 2.730 1.255 ;
        RECT  2.495 0.760 2.615 1.770 ;
        RECT  2.265 0.760 2.495 0.880 ;
        RECT  2.280 1.650 2.495 1.770 ;
        RECT  2.160 1.650 2.280 2.050 ;
        RECT  2.095 0.350 2.265 0.880 ;
        RECT  1.365 1.930 2.160 2.050 ;
        RECT  1.515 0.660 2.095 0.780 ;
        RECT  1.345 0.350 1.515 0.780 ;
        RECT  1.195 1.930 1.365 2.100 ;
    END
END OR4X4AD
MACRO OR4X6AD
    CLASS CORE ;
    FOREIGN OR4X6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.010 0.430 5.200 2.165 ;
        RECT  4.830 0.725 5.010 1.655 ;
        RECT  4.505 0.725 4.830 0.905 ;
        RECT  4.445 1.475 4.830 1.655 ;
        RECT  4.335 0.475 4.505 0.905 ;
        RECT  4.275 1.475 4.445 2.165 ;
        END
        AntennaDiffArea 0.795 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.845 0.880 3.910 1.140 ;
        RECT  3.725 0.880 3.845 1.660 ;
        RECT  1.610 1.540 3.725 1.660 ;
        RECT  1.415 1.290 1.610 1.660 ;
        RECT  1.225 1.290 1.415 1.410 ;
        END
        AntennaGateArea 0.3318 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 0.865 3.570 1.420 ;
        RECT  1.860 1.300 3.430 1.420 ;
        RECT  1.740 1.160 1.860 1.420 ;
        END
        AntennaGateArea 0.331 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.070 0.880 3.190 1.180 ;
        RECT  2.160 1.060 3.070 1.180 ;
        RECT  2.040 0.920 2.160 1.180 ;
        RECT  0.770 0.920 2.040 1.040 ;
        RECT  0.510 0.920 0.770 1.375 ;
        END
        AntennaGateArea 0.331 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.815 2.850 0.935 ;
        RECT  2.330 0.680 2.450 0.935 ;
        RECT  0.320 0.680 2.330 0.800 ;
        RECT  0.200 0.680 0.320 1.430 ;
        RECT  0.070 1.145 0.200 1.375 ;
        END
        AntennaGateArea 0.331 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.865 -0.210 5.320 0.210 ;
        RECT  4.695 -0.210 4.865 0.595 ;
        RECT  4.190 -0.210 4.695 0.210 ;
        RECT  3.930 -0.210 4.190 0.500 ;
        RECT  3.470 -0.210 3.930 0.210 ;
        RECT  3.210 -0.210 3.470 0.500 ;
        RECT  2.730 -0.210 3.210 0.210 ;
        RECT  2.470 -0.210 2.730 0.320 ;
        RECT  1.970 -0.210 2.470 0.210 ;
        RECT  1.710 -0.210 1.970 0.320 ;
        RECT  1.180 -0.210 1.710 0.210 ;
        RECT  0.920 -0.210 1.180 0.560 ;
        RECT  0.000 -0.210 0.920 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.820 2.310 5.320 2.730 ;
        RECT  4.650 1.845 4.820 2.730 ;
        RECT  4.100 2.310 4.650 2.730 ;
        RECT  3.840 2.020 4.100 2.730 ;
        RECT  1.470 2.310 3.840 2.730 ;
        RECT  1.210 2.020 1.470 2.730 ;
        RECT  0.000 2.310 1.210 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.320 2.520 ;
        LAYER M1 ;
        RECT  4.150 1.065 4.585 1.235 ;
        RECT  4.030 0.620 4.150 1.900 ;
        RECT  3.785 0.620 4.030 0.740 ;
        RECT  2.695 1.780 4.030 1.900 ;
        RECT  3.615 0.510 3.785 0.740 ;
        RECT  3.065 0.620 3.615 0.740 ;
        RECT  2.945 0.440 3.065 0.740 ;
        RECT  2.895 0.440 2.945 0.610 ;
        RECT  1.330 0.440 2.895 0.560 ;
        RECT  2.525 1.780 2.695 1.995 ;
        RECT  0.255 1.780 2.525 1.900 ;
        RECT  0.085 1.580 0.255 2.010 ;
    END
END OR4X6AD
MACRO OR4X8AD
    CLASS CORE ;
    FOREIGN OR4X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.325 0.420 6.535 2.145 ;
        RECT  5.850 1.005 6.325 1.605 ;
        RECT  5.680 0.420 5.850 2.190 ;
        RECT  5.625 0.420 5.680 0.850 ;
        RECT  5.650 1.410 5.680 2.190 ;
        END
        AntennaDiffArea 0.844 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.140 0.980 5.260 1.310 ;
        RECT  4.920 1.190 5.140 1.310 ;
        RECT  4.800 1.190 4.920 1.810 ;
        RECT  3.040 1.690 4.800 1.810 ;
        RECT  2.920 1.450 3.040 1.810 ;
        RECT  0.360 1.450 2.920 1.570 ;
        RECT  0.360 0.380 2.185 0.500 ;
        RECT  0.240 0.380 0.360 1.570 ;
        RECT  0.070 0.865 0.240 1.095 ;
        END
        AntennaGateArea 0.438 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.680 0.910 5.015 1.060 ;
        RECT  4.560 0.910 4.680 1.570 ;
        RECT  3.280 1.450 4.560 1.570 ;
        RECT  3.160 1.200 3.280 1.570 ;
        RECT  3.120 1.200 3.160 1.320 ;
        RECT  2.860 1.140 3.120 1.320 ;
        RECT  0.630 1.200 2.860 1.320 ;
        RECT  0.510 0.640 0.630 1.320 ;
        END
        AntennaGateArea 0.438 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.320 0.950 4.440 1.330 ;
        RECT  3.520 1.210 4.320 1.330 ;
        RECT  3.400 0.900 3.520 1.330 ;
        RECT  3.260 0.900 3.400 1.080 ;
        RECT  1.095 0.900 3.260 1.020 ;
        RECT  0.940 0.900 1.095 1.050 ;
        RECT  0.820 0.790 0.940 1.050 ;
        END
        AntennaGateArea 0.438 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.760 0.910 4.160 1.090 ;
        RECT  3.640 0.660 3.760 1.090 ;
        RECT  1.270 0.660 3.640 0.780 ;
        END
        AntennaGateArea 0.438 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.875 -0.210 7.000 0.210 ;
        RECT  6.705 -0.210 6.875 0.815 ;
        RECT  6.155 -0.210 6.705 0.210 ;
        RECT  5.985 -0.210 6.155 0.820 ;
        RECT  5.480 -0.210 5.985 0.210 ;
        RECT  5.220 -0.210 5.480 0.500 ;
        RECT  4.760 -0.210 5.220 0.210 ;
        RECT  4.500 -0.210 4.760 0.500 ;
        RECT  4.020 -0.210 4.500 0.210 ;
        RECT  3.760 -0.210 4.020 0.300 ;
        RECT  3.260 -0.210 3.760 0.210 ;
        RECT  3.000 -0.210 3.260 0.300 ;
        RECT  2.475 -0.210 3.000 0.210 ;
        RECT  2.305 -0.210 2.475 0.525 ;
        RECT  0.000 -0.210 2.305 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.875 2.310 7.000 2.730 ;
        RECT  6.705 1.580 6.875 2.730 ;
        RECT  6.155 2.310 6.705 2.730 ;
        RECT  5.985 1.725 6.155 2.730 ;
        RECT  5.410 2.310 5.985 2.730 ;
        RECT  5.290 1.690 5.410 2.730 ;
        RECT  2.560 2.310 5.290 2.730 ;
        RECT  2.440 1.950 2.560 2.730 ;
        RECT  0.255 2.310 2.440 2.730 ;
        RECT  0.085 1.725 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  5.500 1.000 5.560 1.260 ;
        RECT  5.380 0.635 5.500 1.550 ;
        RECT  5.075 0.635 5.380 0.755 ;
        RECT  5.160 1.430 5.380 1.550 ;
        RECT  5.040 1.430 5.160 2.070 ;
        RECT  4.905 0.470 5.075 0.755 ;
        RECT  2.800 1.950 5.040 2.070 ;
        RECT  4.355 0.635 4.905 0.755 ;
        RECT  4.235 0.420 4.355 0.755 ;
        RECT  4.185 0.420 4.235 0.645 ;
        RECT  2.620 0.420 4.185 0.540 ;
        RECT  2.680 1.705 2.800 2.070 ;
        RECT  1.365 1.705 2.680 1.825 ;
        RECT  1.195 1.705 1.365 2.135 ;
    END
END OR4X8AD
MACRO OR4XLAD
    CLASS CORE ;
    FOREIGN OR4XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 0.690 2.170 1.700 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.000 1.640 1.435 ;
        END
        AntennaGateArea 0.05 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.020 1.330 1.375 ;
        END
        AntennaGateArea 0.05 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.000 0.820 1.465 ;
        END
        AntennaGateArea 0.05 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.000 0.490 1.465 ;
        END
        AntennaGateArea 0.0503 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.765 -0.210 2.240 0.210 ;
        RECT  1.595 -0.210 1.765 0.640 ;
        RECT  0.995 -0.210 1.595 0.210 ;
        RECT  0.825 -0.210 0.995 0.470 ;
        RECT  0.255 -0.210 0.825 0.210 ;
        RECT  0.085 -0.210 0.255 0.640 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.750 2.310 2.240 2.730 ;
        RECT  1.580 1.575 1.750 2.730 ;
        RECT  0.000 2.310 1.580 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.760 0.760 1.880 1.280 ;
        RECT  0.230 0.760 1.760 0.880 ;
        RECT  0.110 0.760 0.230 1.675 ;
    END
END OR4XLAD
MACRO RF1R1WX1AD
    CLASS CORE ;
    FOREIGN RF1R1WX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN WW
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.635 2.010 1.985 2.180 ;
        END
        AntennaGateArea 0.092 ;
    END WW
    PIN WB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.215 1.010 0.240 1.270 ;
        RECT  0.070 1.010 0.215 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END WB
    PIN RWN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 2.005 3.220 2.175 ;
        END
        AntennaGateArea 0.035 ;
    END RWN
    PIN RW
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.910 0.940 3.030 1.255 ;
        RECT  2.905 0.940 2.910 1.060 ;
        RECT  2.785 0.630 2.905 1.060 ;
        RECT  2.545 0.630 2.785 0.770 ;
        END
        AntennaGateArea 0.023 ;
    END RW
    PIN RB
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.200 0.650 3.290 1.655 ;
        RECT  3.150 0.650 3.200 1.860 ;
        RECT  3.055 0.650 3.150 0.820 ;
        RECT  3.060 1.515 3.150 1.860 ;
        END
        AntennaDiffArea 0.135 ;
    END RB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.630 -0.210 3.360 0.210 ;
        RECT  2.370 -0.210 2.630 0.375 ;
        RECT  1.550 -0.210 2.370 0.210 ;
        RECT  1.380 -0.210 1.550 0.395 ;
        RECT  0.240 -0.210 1.380 0.210 ;
        RECT  0.120 -0.210 0.240 0.890 ;
        RECT  0.000 -0.210 0.120 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.605 2.310 3.360 2.730 ;
        RECT  2.435 1.740 2.605 2.730 ;
        RECT  1.515 2.310 2.435 2.730 ;
        RECT  1.345 2.030 1.515 2.730 ;
        RECT  0.230 2.310 1.345 2.730 ;
        RECT  0.110 1.655 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.360 2.520 ;
        LAYER M1 ;
        RECT  2.650 1.180 2.730 1.440 ;
        RECT  2.530 0.960 2.650 1.575 ;
        RECT  2.270 0.960 2.530 1.080 ;
        RECT  2.245 1.455 2.530 1.575 ;
        RECT  1.750 1.210 2.410 1.330 ;
        RECT  2.150 0.625 2.270 1.080 ;
        RECT  2.075 1.455 2.245 1.825 ;
        RECT  1.470 0.960 2.150 1.080 ;
        RECT  1.110 1.680 1.950 1.800 ;
        RECT  1.785 0.550 1.905 0.810 ;
        RECT  1.215 0.550 1.785 0.670 ;
        RECT  1.630 1.210 1.750 1.505 ;
        RECT  0.840 1.385 1.630 1.505 ;
        RECT  1.210 0.960 1.470 1.190 ;
        RECT  1.120 0.380 1.215 0.670 ;
        RECT  1.095 0.330 1.120 0.670 ;
        RECT  0.990 1.680 1.110 2.140 ;
        RECT  0.860 0.330 1.095 0.500 ;
        RECT  0.790 2.020 0.990 2.140 ;
        RECT  0.840 0.630 0.890 0.890 ;
        RECT  0.500 0.380 0.860 0.500 ;
        RECT  0.720 0.630 0.840 1.845 ;
        RECT  0.530 2.020 0.790 2.190 ;
        RECT  0.500 2.020 0.530 2.140 ;
        RECT  0.380 0.380 0.500 2.140 ;
    END
END RF1R1WX1AD
MACRO RF2R1WX1AD
    CLASS CORE ;
    FOREIGN RF2R1WX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN WW
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.635 2.020 1.985 2.190 ;
        END
        AntennaGateArea 0.08 ;
    END WW
    PIN WB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.215 1.010 0.240 1.270 ;
        RECT  0.070 1.010 0.215 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END WB
    PIN R2W
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.110 1.145 5.250 1.375 ;
        RECT  4.960 1.070 5.110 1.440 ;
        END
        AntennaGateArea 0.071 ;
    END R2W
    PIN R2B
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  4.410 0.615 4.495 0.785 ;
        RECT  4.410 1.640 4.495 1.810 ;
        RECT  4.270 0.615 4.410 1.810 ;
        END
        AntennaDiffArea 0.133 ;
    END R2B
    PIN R1W
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.805 1.145 3.850 1.375 ;
        RECT  3.660 0.955 3.805 1.375 ;
        RECT  3.625 0.955 3.660 1.215 ;
        END
        AntennaGateArea 0.071 ;
    END R1W
    PIN R1B
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.035 0.610 3.215 0.780 ;
        RECT  3.035 1.680 3.190 1.945 ;
        RECT  2.915 0.610 3.035 1.945 ;
        RECT  2.870 1.425 2.915 1.945 ;
        END
        AntennaDiffArea 0.133 ;
    END R1B
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.185 -0.210 5.320 0.210 ;
        RECT  5.065 -0.210 5.185 0.895 ;
        RECT  3.910 -0.210 5.065 0.210 ;
        RECT  3.650 -0.210 3.910 0.330 ;
        RECT  2.605 -0.210 3.650 0.210 ;
        RECT  2.435 -0.210 2.605 0.765 ;
        RECT  1.515 -0.210 2.435 0.210 ;
        RECT  1.345 -0.210 1.515 0.460 ;
        RECT  0.240 -0.210 1.345 0.210 ;
        RECT  0.120 -0.210 0.240 0.890 ;
        RECT  0.000 -0.210 0.120 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.185 2.310 5.320 2.730 ;
        RECT  5.065 1.560 5.185 2.730 ;
        RECT  3.845 2.310 5.065 2.730 ;
        RECT  3.675 2.055 3.845 2.730 ;
        RECT  2.605 2.310 3.675 2.730 ;
        RECT  2.435 1.720 2.605 2.730 ;
        RECT  1.515 2.310 2.435 2.730 ;
        RECT  1.345 2.030 1.515 2.730 ;
        RECT  0.230 2.310 1.345 2.730 ;
        RECT  0.110 1.655 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.320 2.520 ;
        LAYER M1 ;
        RECT  4.705 0.635 4.825 1.775 ;
        RECT  4.585 1.205 4.705 1.465 ;
        RECT  3.505 0.625 3.565 0.795 ;
        RECT  3.505 1.560 3.555 1.730 ;
        RECT  3.370 0.625 3.505 1.730 ;
        RECT  3.155 1.165 3.370 1.425 ;
        RECT  2.650 0.960 2.795 1.150 ;
        RECT  2.530 0.960 2.650 1.575 ;
        RECT  2.220 0.960 2.530 1.080 ;
        RECT  2.220 1.455 2.530 1.575 ;
        RECT  1.750 1.210 2.395 1.330 ;
        RECT  2.100 0.580 2.220 1.080 ;
        RECT  2.100 1.455 2.220 1.870 ;
        RECT  1.460 0.960 2.100 1.080 ;
        RECT  1.120 1.655 1.950 1.775 ;
        RECT  1.750 0.580 1.870 0.840 ;
        RECT  1.225 0.580 1.750 0.700 ;
        RECT  1.630 1.210 1.750 1.485 ;
        RECT  0.840 1.365 1.630 1.485 ;
        RECT  1.200 0.960 1.460 1.190 ;
        RECT  1.105 0.380 1.225 0.700 ;
        RECT  1.000 1.655 1.120 2.140 ;
        RECT  1.040 0.380 1.105 0.500 ;
        RECT  0.780 0.330 1.040 0.500 ;
        RECT  0.600 2.020 1.000 2.140 ;
        RECT  0.840 0.630 0.865 0.890 ;
        RECT  0.720 0.630 0.840 1.855 ;
        RECT  0.600 0.380 0.780 0.500 ;
        RECT  0.480 0.380 0.600 2.140 ;
    END
END RF2R1WX1AD
MACRO SDFFHQX1AD
    CLASS CORE ;
    FOREIGN SDFFHQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.560 1.350 3.850 1.655 ;
        END
        AntennaGateArea 0.049 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.080 1.360 3.200 1.620 ;
        RECT  1.890 1.500 3.080 1.620 ;
        RECT  1.770 1.145 1.890 1.620 ;
        RECT  1.520 1.145 1.770 1.415 ;
        END
        AntennaGateArea 0.097 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.910 0.590 8.050 1.810 ;
        RECT  7.850 0.590 7.910 0.850 ;
        RECT  7.850 1.550 7.910 1.810 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.860 2.670 1.120 ;
        END
        AntennaGateArea 0.08 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.930 0.490 1.655 ;
        END
        AntennaGateArea 0.12 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.800 -0.210 8.120 0.210 ;
        RECT  7.540 -0.210 7.800 0.300 ;
        RECT  7.410 -0.210 7.540 0.210 ;
        RECT  7.150 -0.210 7.410 0.300 ;
        RECT  5.845 -0.210 7.150 0.210 ;
        RECT  5.585 -0.210 5.845 0.290 ;
        RECT  3.970 -0.210 5.585 0.210 ;
        RECT  3.710 -0.210 3.970 0.300 ;
        RECT  2.300 -0.210 3.710 0.210 ;
        RECT  2.180 -0.210 2.300 0.500 ;
        RECT  1.110 -0.210 2.180 0.210 ;
        RECT  0.590 -0.210 1.110 0.300 ;
        RECT  0.000 -0.210 0.590 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.700 2.310 8.120 2.730 ;
        RECT  7.440 2.220 7.700 2.730 ;
        RECT  7.290 2.310 7.440 2.730 ;
        RECT  7.030 2.220 7.290 2.730 ;
        RECT  5.835 2.310 7.030 2.730 ;
        RECT  5.575 2.220 5.835 2.730 ;
        RECT  4.650 2.310 5.575 2.730 ;
        RECT  4.390 2.220 4.650 2.730 ;
        RECT  2.580 2.310 4.390 2.730 ;
        RECT  2.320 2.220 2.580 2.730 ;
        RECT  1.940 2.310 2.320 2.730 ;
        RECT  1.680 2.220 1.940 2.730 ;
        RECT  0.570 2.310 1.680 2.730 ;
        RECT  0.350 2.010 0.570 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.120 2.520 ;
        LAYER M1 ;
        RECT  7.525 1.000 7.645 2.100 ;
        RECT  6.950 1.980 7.525 2.100 ;
        RECT  7.340 0.760 7.410 0.880 ;
        RECT  7.220 0.760 7.340 1.590 ;
        RECT  7.150 0.760 7.220 1.260 ;
        RECT  7.035 1.000 7.150 1.260 ;
        RECT  6.830 1.740 6.950 2.100 ;
        RECT  6.745 0.380 6.865 1.580 ;
        RECT  6.435 1.740 6.830 1.860 ;
        RECT  6.575 0.380 6.745 0.500 ;
        RECT  6.555 1.460 6.745 1.580 ;
        RECT  6.505 0.650 6.625 1.050 ;
        RECT  6.315 0.330 6.575 0.500 ;
        RECT  6.435 0.930 6.505 1.050 ;
        RECT  6.245 1.980 6.505 2.190 ;
        RECT  6.315 0.930 6.435 1.860 ;
        RECT  6.195 0.690 6.335 0.810 ;
        RECT  6.110 0.380 6.315 0.500 ;
        RECT  4.940 1.980 6.245 2.100 ;
        RECT  6.075 0.690 6.195 1.860 ;
        RECT  5.990 0.380 6.110 0.540 ;
        RECT  5.965 0.690 6.075 0.890 ;
        RECT  4.630 1.740 6.075 1.860 ;
        RECT  5.420 0.420 5.990 0.540 ;
        RECT  5.855 0.770 5.965 0.890 ;
        RECT  5.835 1.100 5.955 1.360 ;
        RECT  5.595 0.770 5.855 0.960 ;
        RECT  5.465 1.170 5.835 1.290 ;
        RECT  5.345 0.660 5.465 1.620 ;
        RECT  5.300 0.380 5.420 0.540 ;
        RECT  5.180 0.660 5.345 0.780 ;
        RECT  4.855 1.500 5.345 1.620 ;
        RECT  4.900 0.380 5.300 0.500 ;
        RECT  5.050 1.070 5.220 1.325 ;
        RECT  4.860 0.620 5.180 0.780 ;
        RECT  4.150 1.070 5.050 1.190 ;
        RECT  4.770 1.980 4.940 2.190 ;
        RECT  4.640 0.330 4.900 0.500 ;
        RECT  4.500 0.620 4.860 0.740 ;
        RECT  4.300 1.980 4.770 2.100 ;
        RECT  4.260 0.380 4.640 0.500 ;
        RECT  4.510 1.360 4.630 1.860 ;
        RECT  4.345 1.360 4.510 1.480 ;
        RECT  4.180 1.980 4.300 2.140 ;
        RECT  4.140 0.380 4.260 0.540 ;
        RECT  2.835 2.020 4.180 2.140 ;
        RECT  4.090 0.780 4.150 1.615 ;
        RECT  3.620 0.420 4.140 0.540 ;
        RECT  4.030 0.780 4.090 1.900 ;
        RECT  3.390 0.780 4.030 0.900 ;
        RECT  3.970 1.495 4.030 1.900 ;
        RECT  3.560 1.780 3.970 1.900 ;
        RECT  3.440 1.110 3.910 1.230 ;
        RECT  3.500 0.380 3.620 0.540 ;
        RECT  2.540 0.380 3.500 0.500 ;
        RECT  3.320 1.020 3.440 1.860 ;
        RECT  3.270 0.620 3.390 0.900 ;
        RECT  3.150 1.020 3.320 1.140 ;
        RECT  1.650 1.740 3.320 1.860 ;
        RECT  3.070 0.620 3.270 0.740 ;
        RECT  3.030 0.860 3.150 1.140 ;
        RECT  2.910 1.260 2.960 1.380 ;
        RECT  2.910 0.620 2.950 0.740 ;
        RECT  2.790 0.620 2.910 1.380 ;
        RECT  2.715 1.980 2.835 2.140 ;
        RECT  2.690 0.620 2.790 0.740 ;
        RECT  2.700 1.260 2.790 1.380 ;
        RECT  1.150 1.980 2.715 2.100 ;
        RECT  2.420 0.380 2.540 0.740 ;
        RECT  2.150 0.620 2.420 0.740 ;
        RECT  2.150 1.260 2.290 1.380 ;
        RECT  2.030 0.620 2.150 1.380 ;
        RECT  1.730 0.620 2.030 0.785 ;
        RECT  1.140 0.665 1.730 0.785 ;
        RECT  1.610 0.375 1.720 0.495 ;
        RECT  1.530 1.565 1.650 1.860 ;
        RECT  1.390 0.905 1.630 1.025 ;
        RECT  1.460 0.375 1.610 0.540 ;
        RECT  1.390 1.565 1.530 1.685 ;
        RECT  0.230 0.420 1.460 0.540 ;
        RECT  1.270 0.905 1.390 1.685 ;
        RECT  1.030 1.485 1.150 2.100 ;
        RECT  1.020 0.665 1.140 1.270 ;
        RECT  0.730 1.485 1.030 1.605 ;
        RECT  0.850 1.090 1.020 1.270 ;
        RECT  0.780 0.660 0.900 0.920 ;
        RECT  0.730 0.800 0.780 0.920 ;
        RECT  0.610 0.800 0.730 1.605 ;
        RECT  0.110 0.420 0.230 1.745 ;
    END
END SDFFHQX1AD
MACRO SDFFHQX2AD
    CLASS CORE ;
    FOREIGN SDFFHQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 1.350 3.890 1.655 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.070 1.260 3.190 1.660 ;
        RECT  1.890 1.540 3.070 1.660 ;
        RECT  1.770 1.145 1.890 1.660 ;
        RECT  1.540 1.145 1.770 1.415 ;
        END
        AntennaGateArea 0.113 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.730 0.405 8.890 1.930 ;
        END
        AntennaDiffArea 0.363 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.860 2.660 1.160 ;
        END
        AntennaGateArea 0.125 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.145 0.490 1.655 ;
        END
        AntennaGateArea 0.119 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.530 -0.210 8.960 0.210 ;
        RECT  8.270 -0.210 8.530 0.540 ;
        RECT  7.940 -0.210 8.270 0.210 ;
        RECT  7.410 -0.210 7.940 0.300 ;
        RECT  5.800 -0.210 7.410 0.210 ;
        RECT  5.540 -0.210 5.800 0.300 ;
        RECT  4.035 -0.210 5.540 0.210 ;
        RECT  3.775 -0.210 4.035 0.300 ;
        RECT  2.390 -0.210 3.775 0.210 ;
        RECT  2.235 -0.210 2.390 0.500 ;
        RECT  1.220 -0.210 2.235 0.210 ;
        RECT  0.960 -0.210 1.220 0.300 ;
        RECT  0.680 -0.210 0.960 0.210 ;
        RECT  0.420 -0.210 0.680 0.300 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.520 2.310 8.960 2.730 ;
        RECT  8.260 2.220 8.520 2.730 ;
        RECT  8.080 2.310 8.260 2.730 ;
        RECT  7.820 2.220 8.080 2.730 ;
        RECT  7.240 2.310 7.820 2.730 ;
        RECT  6.980 2.220 7.240 2.730 ;
        RECT  5.810 2.310 6.980 2.730 ;
        RECT  5.550 2.210 5.810 2.730 ;
        RECT  4.470 2.310 5.550 2.730 ;
        RECT  4.210 2.260 4.470 2.730 ;
        RECT  2.200 2.310 4.210 2.730 ;
        RECT  1.680 2.260 2.200 2.730 ;
        RECT  0.570 2.310 1.680 2.730 ;
        RECT  0.350 2.020 0.570 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.960 2.520 ;
        LAYER M1 ;
        RECT  8.410 0.980 8.530 2.100 ;
        RECT  7.455 1.980 8.410 2.100 ;
        RECT  8.170 0.760 8.290 1.590 ;
        RECT  7.790 0.760 8.170 0.880 ;
        RECT  8.020 1.330 8.170 1.590 ;
        RECT  7.670 0.760 7.790 1.220 ;
        RECT  7.645 1.000 7.670 1.220 ;
        RECT  7.525 1.405 7.575 1.575 ;
        RECT  7.405 1.110 7.525 1.575 ;
        RECT  7.285 1.715 7.455 2.100 ;
        RECT  7.220 1.110 7.405 1.230 ;
        RECT  7.165 1.470 7.285 2.100 ;
        RECT  7.100 0.420 7.220 1.230 ;
        RECT  6.485 1.470 7.165 1.590 ;
        RECT  6.845 0.420 7.100 0.540 ;
        RECT  6.580 0.720 6.980 0.840 ;
        RECT  6.600 1.715 6.860 1.885 ;
        RECT  6.675 0.355 6.845 0.540 ;
        RECT  5.400 0.420 6.675 0.540 ;
        RECT  6.080 1.715 6.600 1.835 ;
        RECT  6.485 0.720 6.580 1.050 ;
        RECT  6.460 0.720 6.485 1.590 ;
        RECT  6.365 0.930 6.460 1.590 ;
        RECT  6.240 1.470 6.365 1.590 ;
        RECT  6.080 0.670 6.340 0.790 ;
        RECT  6.095 1.955 6.265 2.185 ;
        RECT  4.980 1.955 6.095 2.075 ;
        RECT  5.960 0.670 6.080 1.835 ;
        RECT  5.760 0.670 5.960 0.790 ;
        RECT  5.930 1.500 5.960 1.835 ;
        RECT  4.525 1.715 5.930 1.835 ;
        RECT  5.720 1.090 5.840 1.350 ;
        RECT  5.500 0.670 5.760 0.865 ;
        RECT  5.380 1.180 5.720 1.300 ;
        RECT  5.280 0.380 5.400 0.540 ;
        RECT  5.260 0.660 5.380 1.590 ;
        RECT  4.925 0.380 5.280 0.500 ;
        RECT  5.060 0.660 5.260 0.780 ;
        RECT  4.890 1.470 5.260 1.590 ;
        RECT  4.950 1.070 5.070 1.350 ;
        RECT  4.540 0.620 5.060 0.780 ;
        RECT  4.720 1.955 4.980 2.190 ;
        RECT  4.140 1.070 4.950 1.190 ;
        RECT  4.665 0.330 4.925 0.500 ;
        RECT  1.150 2.020 4.720 2.140 ;
        RECT  4.275 0.380 4.665 0.500 ;
        RECT  4.405 1.385 4.525 1.835 ;
        RECT  4.355 1.385 4.405 1.555 ;
        RECT  4.155 0.380 4.275 0.540 ;
        RECT  3.630 0.420 4.155 0.540 ;
        RECT  4.020 0.780 4.140 1.900 ;
        RECT  3.390 0.780 4.020 0.900 ;
        RECT  3.550 1.780 4.020 1.900 ;
        RECT  3.430 1.110 3.900 1.230 ;
        RECT  3.510 0.380 3.630 0.540 ;
        RECT  2.630 0.380 3.510 0.500 ;
        RECT  3.310 1.020 3.430 1.900 ;
        RECT  3.270 0.620 3.390 0.900 ;
        RECT  3.150 1.020 3.310 1.140 ;
        RECT  1.560 1.780 3.310 1.900 ;
        RECT  3.130 0.620 3.270 0.740 ;
        RECT  3.030 0.880 3.150 1.140 ;
        RECT  2.900 0.620 3.010 0.740 ;
        RECT  2.900 1.300 2.950 1.420 ;
        RECT  2.780 0.620 2.900 1.420 ;
        RECT  2.750 0.620 2.780 0.740 ;
        RECT  2.690 1.300 2.780 1.420 ;
        RECT  2.510 0.380 2.630 0.740 ;
        RECT  2.160 0.620 2.510 0.740 ;
        RECT  2.160 1.300 2.270 1.420 ;
        RECT  2.040 0.620 2.160 1.420 ;
        RECT  1.770 0.620 2.040 0.785 ;
        RECT  2.010 1.300 2.040 1.420 ;
        RECT  1.140 0.665 1.770 0.785 ;
        RECT  1.665 0.360 1.760 0.480 ;
        RECT  1.500 0.360 1.665 0.540 ;
        RECT  1.410 0.905 1.620 1.025 ;
        RECT  1.440 1.575 1.560 1.900 ;
        RECT  0.230 0.420 1.500 0.540 ;
        RECT  1.410 1.575 1.440 1.695 ;
        RECT  1.290 0.905 1.410 1.695 ;
        RECT  1.030 1.495 1.150 2.140 ;
        RECT  1.020 0.665 1.140 1.270 ;
        RECT  0.730 1.495 1.030 1.615 ;
        RECT  0.850 1.090 1.020 1.270 ;
        RECT  0.780 0.660 0.900 0.920 ;
        RECT  0.730 0.800 0.780 0.920 ;
        RECT  0.610 0.800 0.730 1.615 ;
        RECT  0.110 0.420 0.230 1.755 ;
    END
END SDFFHQX2AD
MACRO SDFFHQX4AD
    CLASS CORE ;
    FOREIGN SDFFHQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.690 1.410 4.175 1.610 ;
        END
        AntennaGateArea 0.074 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 0.865 2.450 1.280 ;
        END
        AntennaGateArea 0.15 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.620 1.005 9.730 1.515 ;
        RECT  9.490 0.410 9.620 2.005 ;
        END
        AntennaDiffArea 0.41 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.865 2.930 1.260 ;
        END
        AntennaGateArea 0.112 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.050 1.510 1.220 ;
        RECT  1.075 0.865 1.450 1.220 ;
        END
        AntennaGateArea 0.197 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.995 -0.210 10.080 0.210 ;
        RECT  9.825 -0.210 9.995 0.865 ;
        RECT  9.300 -0.210 9.825 0.210 ;
        RECT  9.040 -0.210 9.300 0.300 ;
        RECT  8.155 -0.210 9.040 0.210 ;
        RECT  7.985 -0.210 8.155 0.255 ;
        RECT  6.575 -0.210 7.985 0.210 ;
        RECT  6.315 -0.210 6.575 0.260 ;
        RECT  4.760 -0.210 6.315 0.210 ;
        RECT  4.500 -0.210 4.760 0.260 ;
        RECT  4.200 -0.210 4.500 0.210 ;
        RECT  3.940 -0.210 4.200 0.260 ;
        RECT  2.520 -0.210 3.940 0.210 ;
        RECT  2.400 -0.210 2.520 0.500 ;
        RECT  1.380 -0.210 2.400 0.210 ;
        RECT  1.120 -0.210 1.380 0.310 ;
        RECT  0.230 -0.210 1.120 0.210 ;
        RECT  0.110 -0.210 0.230 0.860 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.970 2.310 10.080 2.730 ;
        RECT  9.850 1.600 9.970 2.730 ;
        RECT  9.255 2.310 9.850 2.730 ;
        RECT  9.085 2.265 9.255 2.730 ;
        RECT  8.340 2.310 9.085 2.730 ;
        RECT  8.080 2.110 8.340 2.730 ;
        RECT  6.735 2.310 8.080 2.730 ;
        RECT  6.565 2.265 6.735 2.730 ;
        RECT  5.835 2.310 6.565 2.730 ;
        RECT  5.665 2.265 5.835 2.730 ;
        RECT  4.595 2.310 5.665 2.730 ;
        RECT  4.425 2.265 4.595 2.730 ;
        RECT  2.940 2.310 4.425 2.730 ;
        RECT  2.680 2.140 2.940 2.730 ;
        RECT  1.580 2.310 2.680 2.730 ;
        RECT  1.320 2.190 1.580 2.730 ;
        RECT  0.975 2.310 1.320 2.730 ;
        RECT  0.805 1.885 0.975 2.730 ;
        RECT  0.230 2.310 0.805 2.730 ;
        RECT  0.110 1.580 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.080 2.520 ;
        LAYER M1 ;
        RECT  9.250 0.485 9.370 1.980 ;
        RECT  8.830 0.485 9.250 0.605 ;
        RECT  8.990 1.860 9.250 1.980 ;
        RECT  8.730 1.860 8.990 2.070 ;
        RECT  8.795 0.760 8.965 1.740 ;
        RECT  8.570 0.330 8.830 0.605 ;
        RECT  8.300 0.760 8.795 0.880 ;
        RECT  8.270 1.620 8.795 1.740 ;
        RECT  8.130 1.860 8.730 1.980 ;
        RECT  8.060 1.290 8.675 1.410 ;
        RECT  8.180 0.570 8.300 0.880 ;
        RECT  8.010 1.530 8.130 1.980 ;
        RECT  7.940 0.380 8.060 1.410 ;
        RECT  7.555 1.530 8.010 1.650 ;
        RECT  7.230 0.380 7.940 0.500 ;
        RECT  7.770 1.770 7.890 2.030 ;
        RECT  7.040 0.620 7.800 0.740 ;
        RECT  7.195 1.770 7.770 1.895 ;
        RECT  7.525 1.480 7.555 1.650 ;
        RECT  7.385 0.865 7.525 1.650 ;
        RECT  7.350 2.070 7.410 2.190 ;
        RECT  7.160 0.865 7.385 0.985 ;
        RECT  7.150 2.020 7.350 2.190 ;
        RECT  6.970 0.330 7.230 0.500 ;
        RECT  7.040 1.690 7.195 1.895 ;
        RECT  5.040 2.020 7.150 2.140 ;
        RECT  6.920 0.620 7.040 1.895 ;
        RECT  6.160 0.380 6.970 0.500 ;
        RECT  6.710 0.670 6.920 0.790 ;
        RECT  4.670 1.770 6.920 1.895 ;
        RECT  6.490 0.975 6.800 1.235 ;
        RECT  6.455 0.880 6.490 1.235 ;
        RECT  6.335 0.880 6.455 1.650 ;
        RECT  6.040 0.880 6.335 1.000 ;
        RECT  4.975 1.530 6.335 1.650 ;
        RECT  6.080 1.150 6.200 1.410 ;
        RECT  5.900 0.330 6.160 0.500 ;
        RECT  5.370 1.290 6.080 1.410 ;
        RECT  5.920 0.620 6.040 1.000 ;
        RECT  5.260 0.620 5.920 0.740 ;
        RECT  2.760 0.380 5.900 0.500 ;
        RECT  4.910 1.260 5.370 1.410 ;
        RECT  4.780 2.020 5.040 2.190 ;
        RECT  4.790 0.715 4.910 1.410 ;
        RECT  4.415 0.715 4.790 0.835 ;
        RECT  3.350 2.020 4.780 2.140 ;
        RECT  4.550 1.150 4.670 1.895 ;
        RECT  4.295 0.715 4.415 1.860 ;
        RECT  3.570 0.715 4.295 0.835 ;
        RECT  3.980 1.740 4.295 1.860 ;
        RECT  3.885 1.110 4.145 1.255 ;
        RECT  3.720 1.740 3.980 1.900 ;
        RECT  3.570 1.110 3.885 1.230 ;
        RECT  3.310 0.620 3.570 0.835 ;
        RECT  3.450 1.110 3.570 1.760 ;
        RECT  3.410 1.110 3.450 1.260 ;
        RECT  2.930 1.640 3.450 1.760 ;
        RECT  3.290 1.000 3.410 1.260 ;
        RECT  3.230 1.880 3.350 2.140 ;
        RECT  3.170 1.400 3.330 1.520 ;
        RECT  2.690 1.880 3.230 2.000 ;
        RECT  3.050 0.620 3.170 1.520 ;
        RECT  2.900 0.620 3.050 0.740 ;
        RECT  2.810 1.500 2.930 1.760 ;
        RECT  2.505 1.500 2.810 1.620 ;
        RECT  2.640 0.380 2.760 0.740 ;
        RECT  2.570 1.740 2.690 2.000 ;
        RECT  2.280 0.620 2.640 0.740 ;
        RECT  2.165 1.740 2.570 1.860 ;
        RECT  2.335 1.450 2.505 1.620 ;
        RECT  2.140 1.980 2.400 2.190 ;
        RECT  2.040 1.450 2.335 1.570 ;
        RECT  2.160 0.430 2.280 0.740 ;
        RECT  1.995 1.690 2.165 1.860 ;
        RECT  0.615 0.430 2.160 0.550 ;
        RECT  1.820 1.980 2.140 2.100 ;
        RECT  1.920 0.690 2.040 1.570 ;
        RECT  1.750 1.690 1.995 1.810 ;
        RECT  1.700 1.930 1.820 2.100 ;
        RECT  1.630 0.680 1.750 1.810 ;
        RECT  1.260 1.930 1.700 2.050 ;
        RECT  1.570 0.680 1.630 0.940 ;
        RECT  0.955 1.400 1.290 1.520 ;
        RECT  1.140 1.640 1.260 2.050 ;
        RECT  0.615 1.640 1.140 1.760 ;
        RECT  0.835 0.680 0.955 1.520 ;
        RECT  0.785 0.680 0.835 1.260 ;
        RECT  0.620 1.000 0.785 1.260 ;
        RECT  0.475 0.430 0.615 0.810 ;
        RECT  0.475 1.610 0.615 2.040 ;
        RECT  0.445 0.430 0.475 2.040 ;
        RECT  0.350 0.640 0.445 2.040 ;
    END
END SDFFHQX4AD
MACRO SDFFHQX8AD
    CLASS CORE ;
    FOREIGN SDFFHQX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.685 0.940 3.855 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.125 1.205 3.245 1.620 ;
        RECT  1.900 1.500 3.125 1.620 ;
        RECT  1.780 1.145 1.900 1.620 ;
        RECT  1.545 1.145 1.780 1.415 ;
        END
        AntennaGateArea 0.141 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.285 0.420 10.445 2.155 ;
        RECT  9.690 1.005 10.285 1.515 ;
        RECT  9.530 0.420 9.690 2.155 ;
        END
        AntennaDiffArea 0.848 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.860 2.715 1.120 ;
        END
        AntennaGateArea 0.112 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.930 0.490 1.375 ;
        END
        AntennaGateArea 0.201 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.800 -0.210 10.920 0.210 ;
        RECT  10.640 -0.210 10.800 0.875 ;
        RECT  10.080 -0.210 10.640 0.210 ;
        RECT  9.900 -0.210 10.080 0.875 ;
        RECT  9.175 -0.210 9.900 0.210 ;
        RECT  8.650 -0.210 9.175 0.490 ;
        RECT  6.770 -0.210 8.650 0.210 ;
        RECT  6.250 -0.210 6.770 0.265 ;
        RECT  4.355 -0.210 6.250 0.210 ;
        RECT  3.835 -0.210 4.355 0.310 ;
        RECT  2.325 -0.210 3.835 0.210 ;
        RECT  2.160 -0.210 2.325 0.490 ;
        RECT  0.695 -0.210 2.160 0.210 ;
        RECT  0.435 -0.210 0.695 0.310 ;
        RECT  0.000 -0.210 0.435 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.820 2.310 10.920 2.730 ;
        RECT  10.620 1.650 10.820 2.730 ;
        RECT  10.090 2.310 10.620 2.730 ;
        RECT  9.890 1.645 10.090 2.730 ;
        RECT  9.260 2.310 9.890 2.730 ;
        RECT  8.740 2.210 9.260 2.730 ;
        RECT  7.125 2.310 8.740 2.730 ;
        RECT  6.865 2.220 7.125 2.730 ;
        RECT  6.250 2.310 6.865 2.730 ;
        RECT  5.990 2.220 6.250 2.730 ;
        RECT  4.615 2.310 5.990 2.730 ;
        RECT  4.355 2.220 4.615 2.730 ;
        RECT  2.615 2.310 4.355 2.730 ;
        RECT  2.355 2.220 2.615 2.730 ;
        RECT  1.905 2.310 2.355 2.730 ;
        RECT  1.645 2.220 1.905 2.730 ;
        RECT  0.595 2.310 1.645 2.730 ;
        RECT  0.335 2.080 0.595 2.730 ;
        RECT  0.000 2.310 0.335 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.920 2.520 ;
        LAYER M1 ;
        RECT  9.220 1.045 9.410 1.215 ;
        RECT  9.100 1.045 9.220 1.935 ;
        RECT  8.980 1.045 9.100 1.215 ;
        RECT  8.215 1.815 9.100 1.935 ;
        RECT  8.720 1.500 8.980 1.620 ;
        RECT  8.720 0.760 8.940 0.880 ;
        RECT  8.600 0.760 8.720 1.620 ;
        RECT  8.280 0.380 8.400 1.600 ;
        RECT  8.165 0.380 8.280 0.500 ;
        RECT  8.160 1.735 8.215 2.165 ;
        RECT  7.905 0.330 8.165 0.500 ;
        RECT  8.040 0.860 8.160 2.165 ;
        RECT  7.705 0.860 8.040 0.980 ;
        RECT  7.510 1.255 8.040 1.375 ;
        RECT  7.220 0.380 7.905 0.500 ;
        RECT  7.685 1.610 7.855 2.040 ;
        RECT  7.130 1.740 7.685 1.860 ;
        RECT  7.130 0.700 7.585 0.820 ;
        RECT  7.250 1.255 7.510 1.620 ;
        RECT  5.200 1.980 7.350 2.100 ;
        RECT  7.100 0.380 7.220 0.540 ;
        RECT  7.010 0.700 7.130 1.860 ;
        RECT  6.205 0.420 7.100 0.540 ;
        RECT  6.380 0.700 7.010 0.820 ;
        RECT  6.710 1.740 7.010 1.860 ;
        RECT  6.720 1.075 6.890 1.270 ;
        RECT  5.950 1.150 6.720 1.270 ;
        RECT  6.690 1.540 6.710 1.860 ;
        RECT  6.430 1.480 6.690 1.860 ;
        RECT  4.755 1.740 6.430 1.860 ;
        RECT  6.360 0.700 6.380 0.960 ;
        RECT  6.255 0.700 6.360 1.020 ;
        RECT  6.100 0.900 6.255 1.020 ;
        RECT  6.085 0.380 6.205 0.540 ;
        RECT  5.970 0.380 6.085 0.500 ;
        RECT  5.710 0.330 5.970 0.500 ;
        RECT  5.830 0.620 5.950 1.600 ;
        RECT  5.560 0.620 5.830 0.795 ;
        RECT  5.080 1.480 5.830 1.600 ;
        RECT  4.660 0.380 5.710 0.500 ;
        RECT  4.095 0.945 5.700 1.065 ;
        RECT  4.940 0.620 5.560 0.740 ;
        RECT  4.940 1.980 5.200 2.190 ;
        RECT  4.190 1.980 4.940 2.100 ;
        RECT  4.635 1.360 4.755 1.860 ;
        RECT  4.490 0.380 4.660 0.550 ;
        RECT  3.575 0.430 4.490 0.550 ;
        RECT  4.070 1.980 4.190 2.140 ;
        RECT  3.975 0.670 4.095 1.685 ;
        RECT  3.520 2.020 4.070 2.140 ;
        RECT  3.335 0.670 3.975 0.790 ;
        RECT  3.950 1.565 3.975 1.685 ;
        RECT  3.830 1.565 3.950 1.900 ;
        RECT  3.640 1.780 3.830 1.900 ;
        RECT  3.510 1.520 3.710 1.640 ;
        RECT  3.455 0.380 3.575 0.550 ;
        RECT  3.325 1.980 3.520 2.140 ;
        RECT  3.390 0.955 3.510 1.860 ;
        RECT  2.565 0.380 3.455 0.500 ;
        RECT  3.245 0.955 3.390 1.080 ;
        RECT  1.615 1.740 3.390 1.860 ;
        RECT  3.075 0.620 3.335 0.790 ;
        RECT  1.165 1.980 3.325 2.100 ;
        RECT  3.075 0.910 3.245 1.080 ;
        RECT  2.955 1.260 2.995 1.380 ;
        RECT  2.835 0.620 2.955 1.380 ;
        RECT  2.685 0.620 2.835 0.740 ;
        RECT  2.735 1.260 2.835 1.380 ;
        RECT  2.445 0.380 2.565 0.740 ;
        RECT  2.140 0.620 2.445 0.740 ;
        RECT  2.140 1.260 2.325 1.380 ;
        RECT  2.020 0.620 2.140 1.380 ;
        RECT  1.165 0.620 2.020 0.740 ;
        RECT  1.625 0.330 1.745 0.450 ;
        RECT  1.415 0.860 1.655 0.980 ;
        RECT  1.485 0.330 1.625 0.500 ;
        RECT  1.495 1.565 1.615 1.860 ;
        RECT  1.415 1.565 1.495 1.685 ;
        RECT  0.935 0.380 1.485 0.500 ;
        RECT  1.295 0.860 1.415 1.685 ;
        RECT  1.045 0.620 1.165 1.270 ;
        RECT  1.045 1.485 1.165 2.100 ;
        RECT  0.855 1.090 1.045 1.270 ;
        RECT  0.735 1.485 1.045 1.605 ;
        RECT  0.815 0.380 0.935 0.550 ;
        RECT  0.735 0.670 0.915 0.930 ;
        RECT  0.230 0.430 0.815 0.550 ;
        RECT  0.615 0.670 0.735 1.605 ;
        RECT  0.110 0.430 0.230 1.640 ;
    END
END SDFFHQX8AD
MACRO SDFFHX1AD
    CLASS CORE ;
    FOREIGN SDFFHX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.560 1.350 3.850 1.655 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.080 1.360 3.200 1.620 ;
        RECT  1.890 1.500 3.080 1.620 ;
        RECT  1.770 1.145 1.890 1.620 ;
        RECT  1.520 1.145 1.770 1.415 ;
        END
        AntennaGateArea 0.101 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.345 1.740 7.670 1.860 ;
        RECT  7.470 0.690 7.590 0.950 ;
        RECT  7.345 0.830 7.470 0.950 ;
        RECT  7.225 0.830 7.345 1.860 ;
        RECT  7.070 1.425 7.225 1.655 ;
        END
        AntennaDiffArea 0.134 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.190 0.590 8.330 1.810 ;
        RECT  8.130 0.590 8.190 0.850 ;
        RECT  8.130 1.550 8.190 1.810 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.860 2.670 1.120 ;
        END
        AntennaGateArea 0.056 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.930 0.490 1.655 ;
        END
        AntennaGateArea 0.12 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.080 -0.210 8.400 0.210 ;
        RECT  7.820 -0.210 8.080 0.300 ;
        RECT  7.280 -0.210 7.820 0.210 ;
        RECT  7.020 -0.210 7.280 0.300 ;
        RECT  5.845 -0.210 7.020 0.210 ;
        RECT  5.585 -0.210 5.845 0.290 ;
        RECT  3.970 -0.210 5.585 0.210 ;
        RECT  3.710 -0.210 3.970 0.300 ;
        RECT  2.300 -0.210 3.710 0.210 ;
        RECT  2.180 -0.210 2.300 0.500 ;
        RECT  1.110 -0.210 2.180 0.210 ;
        RECT  0.590 -0.210 1.110 0.300 ;
        RECT  0.000 -0.210 0.590 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.980 2.310 8.400 2.730 ;
        RECT  7.720 2.220 7.980 2.730 ;
        RECT  7.290 2.310 7.720 2.730 ;
        RECT  7.030 2.220 7.290 2.730 ;
        RECT  5.835 2.310 7.030 2.730 ;
        RECT  5.575 2.220 5.835 2.730 ;
        RECT  4.650 2.310 5.575 2.730 ;
        RECT  4.390 2.220 4.650 2.730 ;
        RECT  2.580 2.310 4.390 2.730 ;
        RECT  2.320 2.220 2.580 2.730 ;
        RECT  1.940 2.310 2.320 2.730 ;
        RECT  1.680 2.220 1.940 2.730 ;
        RECT  0.570 2.310 1.680 2.730 ;
        RECT  0.350 2.010 0.570 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.400 2.520 ;
        LAYER M1 ;
        RECT  7.950 0.970 8.070 1.430 ;
        RECT  7.925 1.310 7.950 1.430 ;
        RECT  7.805 1.310 7.925 2.100 ;
        RECT  7.710 0.420 7.830 1.190 ;
        RECT  6.950 1.980 7.805 2.100 ;
        RECT  7.105 0.420 7.710 0.540 ;
        RECT  7.620 1.070 7.710 1.190 ;
        RECT  7.500 1.070 7.620 1.590 ;
        RECT  6.985 0.420 7.105 1.260 ;
        RECT  6.830 1.740 6.950 2.100 ;
        RECT  6.745 0.380 6.865 1.580 ;
        RECT  6.435 1.740 6.830 1.860 ;
        RECT  6.575 0.380 6.745 0.500 ;
        RECT  6.555 1.460 6.745 1.580 ;
        RECT  6.505 0.650 6.625 1.050 ;
        RECT  6.315 0.330 6.575 0.500 ;
        RECT  6.435 0.930 6.505 1.050 ;
        RECT  6.245 1.980 6.505 2.190 ;
        RECT  6.315 0.930 6.435 1.860 ;
        RECT  6.195 0.690 6.335 0.810 ;
        RECT  6.110 0.380 6.315 0.500 ;
        RECT  4.940 1.980 6.245 2.100 ;
        RECT  6.075 0.690 6.195 1.860 ;
        RECT  5.990 0.380 6.110 0.540 ;
        RECT  5.965 0.690 6.075 0.890 ;
        RECT  4.630 1.740 6.075 1.860 ;
        RECT  5.420 0.420 5.990 0.540 ;
        RECT  5.855 0.770 5.965 0.890 ;
        RECT  5.835 1.100 5.955 1.360 ;
        RECT  5.595 0.770 5.855 0.960 ;
        RECT  5.465 1.170 5.835 1.290 ;
        RECT  5.345 0.660 5.465 1.620 ;
        RECT  5.300 0.380 5.420 0.540 ;
        RECT  5.180 0.660 5.345 0.780 ;
        RECT  4.855 1.500 5.345 1.620 ;
        RECT  4.900 0.380 5.300 0.500 ;
        RECT  5.050 1.070 5.220 1.325 ;
        RECT  4.860 0.620 5.180 0.780 ;
        RECT  4.150 1.070 5.050 1.190 ;
        RECT  4.770 1.980 4.940 2.190 ;
        RECT  4.640 0.330 4.900 0.500 ;
        RECT  4.500 0.620 4.860 0.740 ;
        RECT  4.300 1.980 4.770 2.100 ;
        RECT  4.260 0.380 4.640 0.500 ;
        RECT  4.510 1.360 4.630 1.860 ;
        RECT  4.345 1.360 4.510 1.480 ;
        RECT  4.180 1.980 4.300 2.140 ;
        RECT  4.140 0.380 4.260 0.540 ;
        RECT  2.835 2.020 4.180 2.140 ;
        RECT  4.090 0.780 4.150 1.615 ;
        RECT  3.620 0.420 4.140 0.540 ;
        RECT  4.030 0.780 4.090 1.900 ;
        RECT  3.390 0.780 4.030 0.900 ;
        RECT  3.970 1.495 4.030 1.900 ;
        RECT  3.560 1.780 3.970 1.900 ;
        RECT  3.440 1.110 3.910 1.230 ;
        RECT  3.500 0.380 3.620 0.540 ;
        RECT  2.540 0.380 3.500 0.500 ;
        RECT  3.320 1.020 3.440 1.860 ;
        RECT  3.270 0.620 3.390 0.900 ;
        RECT  3.150 1.020 3.320 1.140 ;
        RECT  1.650 1.740 3.320 1.860 ;
        RECT  3.070 0.620 3.270 0.740 ;
        RECT  3.030 0.860 3.150 1.140 ;
        RECT  2.910 1.260 2.960 1.380 ;
        RECT  2.910 0.620 2.950 0.740 ;
        RECT  2.790 0.620 2.910 1.380 ;
        RECT  2.715 1.980 2.835 2.140 ;
        RECT  2.690 0.620 2.790 0.740 ;
        RECT  2.700 1.260 2.790 1.380 ;
        RECT  1.150 1.980 2.715 2.100 ;
        RECT  2.420 0.380 2.540 0.740 ;
        RECT  2.150 0.620 2.420 0.740 ;
        RECT  2.150 1.260 2.290 1.380 ;
        RECT  2.030 0.620 2.150 1.380 ;
        RECT  1.730 0.620 2.030 0.785 ;
        RECT  1.140 0.665 1.730 0.785 ;
        RECT  1.610 0.375 1.720 0.495 ;
        RECT  1.530 1.565 1.650 1.860 ;
        RECT  1.390 0.905 1.630 1.025 ;
        RECT  1.460 0.375 1.610 0.540 ;
        RECT  1.390 1.565 1.530 1.685 ;
        RECT  0.230 0.420 1.460 0.540 ;
        RECT  1.270 0.905 1.390 1.685 ;
        RECT  1.030 1.485 1.150 2.100 ;
        RECT  1.020 0.665 1.140 1.270 ;
        RECT  0.730 1.485 1.030 1.605 ;
        RECT  0.850 1.090 1.020 1.270 ;
        RECT  0.780 0.660 0.900 0.920 ;
        RECT  0.730 0.800 0.780 0.920 ;
        RECT  0.610 0.800 0.730 1.605 ;
        RECT  0.110 0.420 0.230 1.745 ;
    END
END SDFFHX1AD
MACRO SDFFHX2AD
    CLASS CORE ;
    FOREIGN SDFFHX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 1.350 3.890 1.655 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.070 1.260 3.190 1.660 ;
        RECT  1.890 1.540 3.070 1.660 ;
        RECT  1.770 1.145 1.890 1.660 ;
        RECT  1.540 1.145 1.770 1.415 ;
        END
        AntennaGateArea 0.117 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.050 1.740 8.460 1.860 ;
        RECT  8.050 0.720 8.330 0.840 ;
        RECT  7.910 0.720 8.050 1.860 ;
        END
        AntennaDiffArea 0.125 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.010 0.405 9.170 1.930 ;
        END
        AntennaDiffArea 0.363 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.860 2.660 1.160 ;
        END
        AntennaGateArea 0.083 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.145 0.490 1.655 ;
        END
        AntennaGateArea 0.12 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.810 -0.210 9.240 0.210 ;
        RECT  8.550 -0.210 8.810 0.300 ;
        RECT  7.940 -0.210 8.550 0.210 ;
        RECT  7.410 -0.210 7.940 0.300 ;
        RECT  5.800 -0.210 7.410 0.210 ;
        RECT  5.540 -0.210 5.800 0.300 ;
        RECT  4.035 -0.210 5.540 0.210 ;
        RECT  3.775 -0.210 4.035 0.300 ;
        RECT  2.390 -0.210 3.775 0.210 ;
        RECT  2.235 -0.210 2.390 0.500 ;
        RECT  1.220 -0.210 2.235 0.210 ;
        RECT  0.960 -0.210 1.220 0.300 ;
        RECT  0.680 -0.210 0.960 0.210 ;
        RECT  0.420 -0.210 0.680 0.300 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.800 2.310 9.240 2.730 ;
        RECT  8.540 2.220 8.800 2.730 ;
        RECT  8.080 2.310 8.540 2.730 ;
        RECT  7.820 2.220 8.080 2.730 ;
        RECT  7.240 2.310 7.820 2.730 ;
        RECT  6.980 2.220 7.240 2.730 ;
        RECT  5.810 2.310 6.980 2.730 ;
        RECT  5.550 2.270 5.810 2.730 ;
        RECT  4.470 2.310 5.550 2.730 ;
        RECT  4.210 2.260 4.470 2.730 ;
        RECT  2.200 2.310 4.210 2.730 ;
        RECT  1.680 2.260 2.200 2.730 ;
        RECT  0.570 2.310 1.680 2.730 ;
        RECT  0.350 2.020 0.570 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.240 2.520 ;
        LAYER M1 ;
        RECT  8.690 0.980 8.810 2.100 ;
        RECT  7.455 1.980 8.690 2.100 ;
        RECT  8.450 0.420 8.570 1.590 ;
        RECT  8.420 0.420 8.450 0.540 ;
        RECT  8.300 1.330 8.450 1.590 ;
        RECT  8.160 0.380 8.420 0.540 ;
        RECT  7.790 0.420 8.160 0.540 ;
        RECT  7.670 0.420 7.790 1.220 ;
        RECT  7.645 1.000 7.670 1.220 ;
        RECT  7.525 1.405 7.575 1.575 ;
        RECT  7.405 1.110 7.525 1.575 ;
        RECT  7.285 1.715 7.455 2.100 ;
        RECT  7.220 1.110 7.405 1.230 ;
        RECT  7.165 1.470 7.285 2.100 ;
        RECT  7.100 0.420 7.220 1.230 ;
        RECT  6.485 1.470 7.165 1.590 ;
        RECT  6.845 0.420 7.100 0.540 ;
        RECT  6.580 0.720 6.980 0.840 ;
        RECT  6.600 1.715 6.860 1.895 ;
        RECT  6.675 0.355 6.845 0.540 ;
        RECT  5.290 0.420 6.675 0.540 ;
        RECT  6.080 1.715 6.600 1.835 ;
        RECT  6.485 0.720 6.580 1.050 ;
        RECT  6.460 0.720 6.485 1.590 ;
        RECT  6.365 0.930 6.460 1.590 ;
        RECT  6.240 1.470 6.365 1.590 ;
        RECT  6.080 0.670 6.340 0.790 ;
        RECT  6.095 1.955 6.265 2.185 ;
        RECT  4.980 1.955 6.095 2.075 ;
        RECT  5.960 0.670 6.080 1.835 ;
        RECT  5.760 0.670 5.960 0.790 ;
        RECT  5.930 1.500 5.960 1.835 ;
        RECT  4.525 1.715 5.930 1.835 ;
        RECT  5.720 1.090 5.840 1.350 ;
        RECT  5.500 0.670 5.760 0.865 ;
        RECT  5.380 1.180 5.720 1.300 ;
        RECT  5.260 0.660 5.380 1.590 ;
        RECT  5.170 0.380 5.290 0.540 ;
        RECT  5.050 0.660 5.260 0.780 ;
        RECT  4.890 1.470 5.260 1.590 ;
        RECT  4.925 0.380 5.170 0.500 ;
        RECT  4.950 1.070 5.070 1.350 ;
        RECT  4.530 0.620 5.050 0.780 ;
        RECT  4.720 1.955 4.980 2.190 ;
        RECT  4.140 1.070 4.950 1.190 ;
        RECT  4.665 0.330 4.925 0.500 ;
        RECT  1.150 2.020 4.720 2.140 ;
        RECT  4.275 0.380 4.665 0.500 ;
        RECT  4.405 1.385 4.525 1.835 ;
        RECT  4.355 1.385 4.405 1.555 ;
        RECT  4.155 0.380 4.275 0.540 ;
        RECT  3.630 0.420 4.155 0.540 ;
        RECT  4.020 0.780 4.140 1.900 ;
        RECT  3.390 0.780 4.020 0.900 ;
        RECT  3.550 1.780 4.020 1.900 ;
        RECT  3.430 1.110 3.900 1.230 ;
        RECT  3.510 0.380 3.630 0.540 ;
        RECT  2.630 0.380 3.510 0.500 ;
        RECT  3.310 1.020 3.430 1.900 ;
        RECT  3.270 0.620 3.390 0.900 ;
        RECT  3.150 1.020 3.310 1.140 ;
        RECT  1.560 1.780 3.310 1.900 ;
        RECT  3.130 0.620 3.270 0.740 ;
        RECT  3.030 0.880 3.150 1.140 ;
        RECT  2.900 0.620 3.010 0.740 ;
        RECT  2.900 1.300 2.950 1.420 ;
        RECT  2.780 0.620 2.900 1.420 ;
        RECT  2.750 0.620 2.780 0.740 ;
        RECT  2.690 1.300 2.780 1.420 ;
        RECT  2.510 0.380 2.630 0.740 ;
        RECT  2.160 0.620 2.510 0.740 ;
        RECT  2.160 1.300 2.270 1.420 ;
        RECT  2.040 0.620 2.160 1.420 ;
        RECT  1.770 0.620 2.040 0.785 ;
        RECT  2.010 1.300 2.040 1.420 ;
        RECT  1.140 0.665 1.770 0.785 ;
        RECT  1.665 0.380 1.760 0.500 ;
        RECT  1.500 0.380 1.665 0.540 ;
        RECT  1.410 0.905 1.620 1.025 ;
        RECT  1.440 1.575 1.560 1.900 ;
        RECT  0.230 0.420 1.500 0.540 ;
        RECT  1.410 1.575 1.440 1.695 ;
        RECT  1.290 0.905 1.410 1.695 ;
        RECT  1.030 1.495 1.150 2.140 ;
        RECT  1.020 0.665 1.140 1.270 ;
        RECT  0.730 1.495 1.030 1.615 ;
        RECT  0.850 1.090 1.020 1.270 ;
        RECT  0.780 0.660 0.900 0.920 ;
        RECT  0.730 0.800 0.780 0.920 ;
        RECT  0.610 0.800 0.730 1.615 ;
        RECT  0.110 0.420 0.230 1.755 ;
    END
END SDFFHX2AD
MACRO SDFFHX4AD
    CLASS CORE ;
    FOREIGN SDFFHX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.690 1.410 4.175 1.610 ;
        END
        AntennaGateArea 0.074 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 0.865 2.450 1.280 ;
        END
        AntennaGateArea 0.15 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.235 1.750 9.635 1.890 ;
        RECT  9.235 0.760 9.450 0.890 ;
        RECT  9.105 0.760 9.235 1.890 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.180 1.005 10.290 1.515 ;
        RECT  10.050 0.410 10.180 2.005 ;
        END
        AntennaDiffArea 0.41 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.865 2.930 1.260 ;
        END
        AntennaGateArea 0.112 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.450 1.050 1.510 1.220 ;
        RECT  1.075 0.865 1.450 1.220 ;
        END
        AntennaGateArea 0.197 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.555 -0.210 10.640 0.210 ;
        RECT  10.385 -0.210 10.555 0.865 ;
        RECT  9.860 -0.210 10.385 0.210 ;
        RECT  9.600 -0.210 9.860 0.300 ;
        RECT  9.060 -0.210 9.600 0.210 ;
        RECT  8.800 -0.210 9.060 0.300 ;
        RECT  8.475 -0.210 8.800 0.210 ;
        RECT  8.215 -0.210 8.475 0.300 ;
        RECT  6.670 -0.210 8.215 0.210 ;
        RECT  6.410 -0.210 6.670 0.260 ;
        RECT  4.760 -0.210 6.410 0.210 ;
        RECT  4.500 -0.210 4.760 0.260 ;
        RECT  4.200 -0.210 4.500 0.210 ;
        RECT  3.940 -0.210 4.200 0.260 ;
        RECT  2.520 -0.210 3.940 0.210 ;
        RECT  2.400 -0.210 2.520 0.500 ;
        RECT  1.380 -0.210 2.400 0.210 ;
        RECT  1.120 -0.210 1.380 0.310 ;
        RECT  0.230 -0.210 1.120 0.210 ;
        RECT  0.110 -0.210 0.230 0.860 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.530 2.310 10.640 2.730 ;
        RECT  10.410 1.600 10.530 2.730 ;
        RECT  9.815 2.310 10.410 2.730 ;
        RECT  9.645 2.265 9.815 2.730 ;
        RECT  9.125 2.310 9.645 2.730 ;
        RECT  8.955 2.265 9.125 2.730 ;
        RECT  8.375 2.310 8.955 2.730 ;
        RECT  8.115 2.220 8.375 2.730 ;
        RECT  6.735 2.310 8.115 2.730 ;
        RECT  6.565 2.265 6.735 2.730 ;
        RECT  5.835 2.310 6.565 2.730 ;
        RECT  5.665 2.265 5.835 2.730 ;
        RECT  4.595 2.310 5.665 2.730 ;
        RECT  4.425 2.265 4.595 2.730 ;
        RECT  2.940 2.310 4.425 2.730 ;
        RECT  2.680 2.140 2.940 2.730 ;
        RECT  1.580 2.310 2.680 2.730 ;
        RECT  1.320 2.190 1.580 2.730 ;
        RECT  0.975 2.310 1.320 2.730 ;
        RECT  0.805 1.885 0.975 2.730 ;
        RECT  0.230 2.310 0.805 2.730 ;
        RECT  0.110 1.580 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.640 2.520 ;
        LAYER M1 ;
        RECT  9.810 0.990 9.930 2.140 ;
        RECT  8.910 2.020 9.810 2.140 ;
        RECT  9.570 0.420 9.690 1.545 ;
        RECT  8.970 0.420 9.570 0.540 ;
        RECT  9.355 1.375 9.570 1.545 ;
        RECT  8.850 0.420 8.970 1.230 ;
        RECT  8.790 1.750 8.910 2.140 ;
        RECT  8.820 0.970 8.850 1.230 ;
        RECT  8.450 1.750 8.790 1.870 ;
        RECT  8.570 0.420 8.690 1.620 ;
        RECT  8.095 0.420 8.570 0.540 ;
        RECT  8.330 0.690 8.450 1.870 ;
        RECT  7.550 1.480 8.330 1.600 ;
        RECT  7.975 0.380 8.095 0.540 ;
        RECT  7.305 0.380 7.975 0.500 ;
        RECT  7.740 1.770 7.910 1.950 ;
        RECT  7.105 0.620 7.875 0.740 ;
        RECT  7.225 1.770 7.740 1.895 ;
        RECT  7.485 1.480 7.550 1.650 ;
        RECT  7.345 0.865 7.485 1.650 ;
        RECT  7.145 2.020 7.405 2.190 ;
        RECT  7.225 0.865 7.345 0.985 ;
        RECT  7.045 0.330 7.305 0.500 ;
        RECT  7.105 1.690 7.225 1.895 ;
        RECT  5.040 2.020 7.145 2.140 ;
        RECT  6.985 0.620 7.105 1.895 ;
        RECT  6.160 0.380 7.045 0.500 ;
        RECT  6.805 0.670 6.985 0.790 ;
        RECT  6.695 1.770 6.985 1.895 ;
        RECT  6.490 0.950 6.850 1.070 ;
        RECT  6.575 1.215 6.695 1.895 ;
        RECT  4.670 1.770 6.575 1.895 ;
        RECT  6.455 0.880 6.490 1.070 ;
        RECT  6.335 0.880 6.455 1.650 ;
        RECT  6.040 0.880 6.335 1.000 ;
        RECT  4.975 1.530 6.335 1.650 ;
        RECT  6.080 1.150 6.200 1.410 ;
        RECT  5.900 0.330 6.160 0.500 ;
        RECT  5.370 1.290 6.080 1.410 ;
        RECT  5.920 0.620 6.040 1.000 ;
        RECT  5.260 0.620 5.920 0.740 ;
        RECT  2.760 0.380 5.900 0.500 ;
        RECT  4.910 1.260 5.370 1.410 ;
        RECT  4.780 2.020 5.040 2.190 ;
        RECT  4.790 0.715 4.910 1.410 ;
        RECT  4.415 0.715 4.790 0.835 ;
        RECT  3.350 2.020 4.780 2.140 ;
        RECT  4.550 1.150 4.670 1.895 ;
        RECT  4.295 0.715 4.415 1.860 ;
        RECT  3.570 0.715 4.295 0.835 ;
        RECT  3.980 1.740 4.295 1.860 ;
        RECT  3.885 1.110 4.145 1.255 ;
        RECT  3.720 1.740 3.980 1.900 ;
        RECT  3.570 1.110 3.885 1.230 ;
        RECT  3.310 0.620 3.570 0.835 ;
        RECT  3.450 1.110 3.570 1.760 ;
        RECT  3.410 1.110 3.450 1.260 ;
        RECT  2.930 1.640 3.450 1.760 ;
        RECT  3.290 1.000 3.410 1.260 ;
        RECT  3.230 1.880 3.350 2.140 ;
        RECT  3.170 1.400 3.330 1.520 ;
        RECT  2.690 1.880 3.230 2.000 ;
        RECT  3.050 0.620 3.170 1.520 ;
        RECT  2.900 0.620 3.050 0.740 ;
        RECT  2.810 1.500 2.930 1.760 ;
        RECT  2.505 1.500 2.810 1.620 ;
        RECT  2.640 0.380 2.760 0.740 ;
        RECT  2.570 1.740 2.690 2.000 ;
        RECT  2.280 0.620 2.640 0.740 ;
        RECT  2.165 1.740 2.570 1.860 ;
        RECT  2.335 1.450 2.505 1.620 ;
        RECT  2.140 1.980 2.400 2.190 ;
        RECT  2.040 1.450 2.335 1.570 ;
        RECT  2.160 0.430 2.280 0.740 ;
        RECT  1.995 1.690 2.165 1.860 ;
        RECT  0.615 0.430 2.160 0.550 ;
        RECT  1.820 1.980 2.140 2.100 ;
        RECT  1.920 0.690 2.040 1.570 ;
        RECT  1.750 1.690 1.995 1.810 ;
        RECT  1.700 1.930 1.820 2.100 ;
        RECT  1.630 0.680 1.750 1.810 ;
        RECT  1.260 1.930 1.700 2.050 ;
        RECT  1.570 0.680 1.630 0.940 ;
        RECT  0.955 1.400 1.290 1.520 ;
        RECT  1.140 1.640 1.260 2.050 ;
        RECT  0.615 1.640 1.140 1.760 ;
        RECT  0.835 0.680 0.955 1.520 ;
        RECT  0.785 0.680 0.835 1.260 ;
        RECT  0.620 1.000 0.785 1.260 ;
        RECT  0.475 0.430 0.615 0.810 ;
        RECT  0.475 1.610 0.615 2.040 ;
        RECT  0.445 0.430 0.475 2.040 ;
        RECT  0.350 0.640 0.445 2.040 ;
    END
END SDFFHX4AD
MACRO SDFFHX8AD
    CLASS CORE ;
    FOREIGN SDFFHX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.160 1.300 7.535 1.610 ;
        END
        AntennaGateArea 0.139 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.570 0.865 3.740 0.990 ;
        RECT  3.240 0.865 3.570 1.095 ;
        END
        AntennaGateArea 0.269 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.100 1.710 16.335 1.900 ;
        RECT  15.930 0.640 16.100 1.900 ;
        RECT  15.900 0.640 15.930 0.900 ;
        RECT  15.610 1.285 15.930 1.795 ;
        END
        AntennaDiffArea 0.124 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  17.570 0.410 17.770 2.005 ;
        RECT  17.035 1.005 17.570 1.515 ;
        RECT  16.865 0.410 17.035 2.005 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.910 1.105 4.430 1.255 ;
        RECT  3.850 1.135 3.910 1.255 ;
        RECT  3.710 1.135 3.850 1.375 ;
        END
        AntennaGateArea 0.279 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.065 1.770 1.235 ;
        RECT  1.340 0.865 1.720 1.235 ;
        END
        AntennaGateArea 0.353 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.115 -0.210 18.200 0.210 ;
        RECT  17.945 -0.210 18.115 0.865 ;
        RECT  17.395 -0.210 17.945 0.210 ;
        RECT  17.225 -0.210 17.395 0.865 ;
        RECT  16.605 -0.210 17.225 0.210 ;
        RECT  16.435 -0.210 16.605 0.260 ;
        RECT  15.680 -0.210 16.435 0.210 ;
        RECT  15.510 -0.210 15.680 0.260 ;
        RECT  12.720 -0.210 15.510 0.210 ;
        RECT  12.550 -0.210 12.720 0.260 ;
        RECT  11.960 -0.210 12.550 0.210 ;
        RECT  11.790 -0.210 11.960 0.260 ;
        RECT  11.200 -0.210 11.790 0.210 ;
        RECT  11.030 -0.210 11.200 0.260 ;
        RECT  9.900 -0.210 11.030 0.210 ;
        RECT  9.640 -0.210 9.900 0.430 ;
        RECT  8.460 -0.210 9.640 0.210 ;
        RECT  8.290 -0.210 8.460 0.260 ;
        RECT  7.090 -0.210 8.290 0.210 ;
        RECT  6.970 -0.210 7.090 0.450 ;
        RECT  4.700 -0.210 6.970 0.210 ;
        RECT  4.580 -0.210 4.700 0.500 ;
        RECT  3.475 -0.210 4.580 0.210 ;
        RECT  2.780 -0.210 3.475 0.455 ;
        RECT  1.670 -0.210 2.780 0.210 ;
        RECT  1.410 -0.210 1.670 0.310 ;
        RECT  0.590 -0.210 1.410 0.210 ;
        RECT  0.470 -0.210 0.590 0.860 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  18.115 2.310 18.200 2.730 ;
        RECT  17.945 1.645 18.115 2.730 ;
        RECT  17.395 2.310 17.945 2.730 ;
        RECT  17.225 1.725 17.395 2.730 ;
        RECT  16.605 2.310 17.225 2.730 ;
        RECT  16.435 2.260 16.605 2.730 ;
        RECT  15.910 2.310 16.435 2.730 ;
        RECT  15.740 2.260 15.910 2.730 ;
        RECT  12.530 2.310 15.740 2.730 ;
        RECT  12.360 2.220 12.530 2.730 ;
        RECT  11.770 2.310 12.360 2.730 ;
        RECT  11.600 2.220 11.770 2.730 ;
        RECT  11.035 2.310 11.600 2.730 ;
        RECT  10.865 2.220 11.035 2.730 ;
        RECT  9.615 2.310 10.865 2.730 ;
        RECT  9.445 2.220 9.615 2.730 ;
        RECT  8.240 2.310 9.445 2.730 ;
        RECT  7.980 2.220 8.240 2.730 ;
        RECT  4.770 2.310 7.980 2.730 ;
        RECT  4.510 2.105 4.770 2.730 ;
        RECT  4.370 2.310 4.510 2.730 ;
        RECT  4.110 2.105 4.370 2.730 ;
        RECT  3.670 2.310 4.110 2.730 ;
        RECT  3.410 2.105 3.670 2.730 ;
        RECT  2.030 2.310 3.410 2.730 ;
        RECT  1.770 2.190 2.030 2.730 ;
        RECT  1.380 2.310 1.770 2.730 ;
        RECT  1.120 2.040 1.380 2.730 ;
        RECT  0.590 2.310 1.120 2.730 ;
        RECT  0.470 1.575 0.590 2.730 ;
        RECT  0.000 2.310 0.470 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 18.200 2.520 ;
        LAYER M1 ;
        RECT  16.610 1.035 16.730 2.140 ;
        RECT  16.560 1.035 16.610 1.205 ;
        RECT  15.410 2.020 16.610 2.140 ;
        RECT  16.290 0.380 16.410 1.590 ;
        RECT  16.270 0.380 16.290 0.500 ;
        RECT  16.220 1.330 16.290 1.590 ;
        RECT  16.010 0.350 16.270 0.500 ;
        RECT  15.780 0.380 16.010 0.500 ;
        RECT  15.660 0.380 15.780 1.165 ;
        RECT  15.610 0.995 15.660 1.165 ;
        RECT  15.370 0.380 15.490 1.725 ;
        RECT  15.290 1.845 15.410 2.140 ;
        RECT  13.010 0.380 15.370 0.500 ;
        RECT  15.210 1.845 15.290 1.965 ;
        RECT  15.090 0.640 15.210 1.965 ;
        RECT  14.995 0.640 15.090 0.985 ;
        RECT  13.435 1.505 15.090 1.625 ;
        RECT  13.420 0.865 14.995 0.985 ;
        RECT  12.280 0.620 14.845 0.740 ;
        RECT  13.385 1.785 14.780 1.905 ;
        RECT  13.285 1.740 13.385 1.905 ;
        RECT  12.280 1.740 13.285 1.860 ;
        RECT  12.885 1.980 13.145 2.145 ;
        RECT  12.840 0.330 13.010 0.500 ;
        RECT  8.800 1.980 12.885 2.100 ;
        RECT  10.145 0.380 12.840 0.500 ;
        RECT  12.160 0.620 12.280 1.860 ;
        RECT  11.365 0.620 12.160 0.740 ;
        RECT  11.435 1.740 12.160 1.860 ;
        RECT  10.760 0.950 12.025 1.070 ;
        RECT  11.175 1.400 11.435 1.860 ;
        RECT  10.960 1.660 11.175 1.860 ;
        RECT  8.400 1.740 10.960 1.860 ;
        RECT  10.640 0.690 10.760 1.620 ;
        RECT  10.445 0.690 10.640 0.910 ;
        RECT  8.730 1.500 10.640 1.620 ;
        RECT  9.070 1.030 10.520 1.190 ;
        RECT  9.240 0.790 10.445 0.910 ;
        RECT  10.025 0.380 10.145 0.670 ;
        RECT  9.480 0.550 10.025 0.670 ;
        RECT  9.360 0.380 9.480 0.670 ;
        RECT  7.330 0.380 9.360 0.500 ;
        RECT  9.170 0.780 9.240 0.910 ;
        RECT  8.910 0.740 9.170 0.910 ;
        RECT  8.950 1.030 9.070 1.290 ;
        RECT  8.160 1.030 8.950 1.150 ;
        RECT  8.540 1.980 8.800 2.190 ;
        RECT  7.710 1.980 8.540 2.100 ;
        RECT  8.280 1.300 8.400 1.860 ;
        RECT  8.040 0.745 8.160 1.860 ;
        RECT  7.790 0.745 8.040 0.865 ;
        RECT  7.470 1.740 8.040 1.860 ;
        RECT  7.800 1.060 7.920 1.365 ;
        RECT  7.010 1.060 7.800 1.180 ;
        RECT  7.530 0.620 7.790 0.940 ;
        RECT  7.590 1.980 7.710 2.140 ;
        RECT  5.430 2.020 7.590 2.140 ;
        RECT  6.610 0.820 7.530 0.940 ;
        RECT  7.280 1.740 7.470 1.900 ;
        RECT  7.210 0.380 7.330 0.690 ;
        RECT  6.080 1.780 7.280 1.900 ;
        RECT  6.850 0.570 7.210 0.690 ;
        RECT  6.890 1.060 7.010 1.660 ;
        RECT  6.370 1.060 6.890 1.180 ;
        RECT  5.430 1.540 6.890 1.660 ;
        RECT  6.730 0.380 6.850 0.690 ;
        RECT  6.130 1.300 6.770 1.420 ;
        RECT  4.940 0.380 6.730 0.500 ;
        RECT  6.490 0.620 6.610 0.940 ;
        RECT  6.300 0.620 6.490 0.780 ;
        RECT  6.250 0.920 6.370 1.180 ;
        RECT  5.490 0.620 6.300 0.740 ;
        RECT  5.900 0.860 6.130 1.420 ;
        RECT  5.235 0.860 5.900 0.980 ;
        RECT  5.150 1.300 5.900 1.420 ;
        RECT  5.310 1.540 5.430 1.745 ;
        RECT  5.310 1.865 5.430 2.140 ;
        RECT  4.005 1.625 5.310 1.745 ;
        RECT  3.165 1.865 5.310 1.985 ;
        RECT  5.115 0.630 5.235 0.980 ;
        RECT  4.890 1.300 5.150 1.505 ;
        RECT  4.220 0.860 5.115 0.980 ;
        RECT  4.820 0.380 4.940 0.740 ;
        RECT  4.130 1.385 4.890 1.505 ;
        RECT  4.460 0.620 4.820 0.740 ;
        RECT  4.340 0.380 4.460 0.740 ;
        RECT  3.980 0.380 4.340 0.500 ;
        RECT  4.100 0.620 4.220 0.980 ;
        RECT  3.835 1.540 4.005 1.745 ;
        RECT  3.860 0.380 3.980 0.745 ;
        RECT  2.560 0.625 3.860 0.745 ;
        RECT  3.425 1.540 3.835 1.660 ;
        RECT  3.305 1.430 3.425 1.660 ;
        RECT  2.320 1.430 3.305 1.550 ;
        RECT  3.045 1.740 3.165 1.985 ;
        RECT  2.965 1.740 3.045 1.860 ;
        RECT  2.445 1.690 2.965 1.860 ;
        RECT  2.590 1.980 2.850 2.190 ;
        RECT  2.270 1.980 2.590 2.100 ;
        RECT  2.440 0.430 2.560 0.745 ;
        RECT  2.050 1.690 2.445 1.810 ;
        RECT  1.020 0.430 2.440 0.550 ;
        RECT  2.200 0.675 2.320 1.550 ;
        RECT  2.150 1.930 2.270 2.100 ;
        RECT  1.620 1.930 2.150 2.050 ;
        RECT  1.930 0.670 2.050 1.810 ;
        RECT  1.860 0.670 1.930 0.930 ;
        RECT  1.220 1.500 1.650 1.660 ;
        RECT  1.500 1.800 1.620 2.050 ;
        RECT  0.975 1.800 1.500 1.920 ;
        RECT  1.100 0.690 1.220 1.660 ;
        RECT  0.980 1.000 1.100 1.260 ;
        RECT  0.835 0.400 1.020 0.550 ;
        RECT  0.835 1.620 0.975 2.050 ;
        RECT  0.710 0.400 0.835 2.050 ;
        RECT  0.230 1.145 0.710 1.265 ;
        RECT  0.110 0.510 0.230 2.095 ;
    END
END SDFFHX8AD
MACRO SDFFNHX1AD
    CLASS CORE ;
    FOREIGN SDFFNHX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.320 1.350 3.570 1.655 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 2.030 2.215 2.190 ;
        END
        AntennaGateArea 0.096 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.170 0.680 7.290 0.940 ;
        RECT  7.030 0.760 7.170 0.940 ;
        RECT  7.030 1.730 7.145 1.850 ;
        RECT  6.910 0.760 7.030 1.850 ;
        RECT  6.790 1.425 6.910 1.850 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.010 1.145 8.050 1.375 ;
        RECT  7.890 0.610 8.010 1.910 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.980 2.570 1.240 ;
        RECT  2.305 0.860 2.450 1.350 ;
        END
        AntennaGateArea 0.061 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.125 1.330 1.375 ;
        RECT  1.020 1.025 1.190 1.375 ;
        END
        AntennaGateArea 0.118 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.815 -0.210 8.120 0.210 ;
        RECT  7.645 -0.210 7.815 0.360 ;
        RECT  6.970 -0.210 7.645 0.210 ;
        RECT  6.710 -0.210 6.970 0.300 ;
        RECT  5.600 -0.210 6.710 0.210 ;
        RECT  5.340 -0.210 5.600 0.300 ;
        RECT  3.855 -0.210 5.340 0.210 ;
        RECT  3.595 -0.210 3.855 0.310 ;
        RECT  2.170 -0.210 3.595 0.210 ;
        RECT  1.910 -0.210 2.170 0.380 ;
        RECT  1.265 -0.210 1.910 0.210 ;
        RECT  1.095 -0.210 1.265 0.375 ;
        RECT  0.335 -0.210 1.095 0.210 ;
        RECT  0.165 -0.210 0.335 0.405 ;
        RECT  0.000 -0.210 0.165 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.630 2.310 8.120 2.730 ;
        RECT  7.510 1.885 7.630 2.730 ;
        RECT  6.755 2.310 7.510 2.730 ;
        RECT  6.495 2.220 6.755 2.730 ;
        RECT  5.395 2.310 6.495 2.730 ;
        RECT  5.135 2.220 5.395 2.730 ;
        RECT  4.365 2.310 5.135 2.730 ;
        RECT  4.105 2.220 4.365 2.730 ;
        RECT  2.595 2.310 4.105 2.730 ;
        RECT  2.335 2.070 2.595 2.730 ;
        RECT  1.220 2.310 2.335 2.730 ;
        RECT  0.960 1.965 1.220 2.730 ;
        RECT  0.255 2.310 0.960 2.730 ;
        RECT  0.085 1.540 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.120 2.520 ;
        LAYER M1 ;
        RECT  7.650 1.000 7.770 1.760 ;
        RECT  7.390 1.640 7.650 1.760 ;
        RECT  7.410 0.405 7.530 1.520 ;
        RECT  7.150 0.405 7.410 0.555 ;
        RECT  7.150 1.400 7.410 1.520 ;
        RECT  7.270 1.640 7.390 2.100 ;
        RECT  6.310 1.980 7.270 2.100 ;
        RECT  6.770 0.435 7.150 0.555 ;
        RECT  6.650 0.435 6.770 1.270 ;
        RECT  6.410 0.380 6.530 1.550 ;
        RECT  6.240 0.380 6.410 0.500 ;
        RECT  6.255 1.430 6.410 1.550 ;
        RECT  6.190 1.810 6.310 2.100 ;
        RECT  6.170 0.680 6.290 1.050 ;
        RECT  6.135 1.430 6.255 1.690 ;
        RECT  5.980 0.330 6.240 0.500 ;
        RECT  6.015 1.810 6.190 1.930 ;
        RECT  6.015 0.930 6.170 1.050 ;
        RECT  5.895 0.930 6.015 1.930 ;
        RECT  5.775 0.660 6.000 0.780 ;
        RECT  5.855 0.380 5.980 0.500 ;
        RECT  5.715 2.070 5.965 2.190 ;
        RECT  5.735 0.380 5.855 0.540 ;
        RECT  5.655 0.660 5.775 1.860 ;
        RECT  5.130 0.420 5.735 0.540 ;
        RECT  5.595 1.980 5.715 2.190 ;
        RECT  5.160 0.660 5.655 0.780 ;
        RECT  4.270 1.740 5.655 1.860 ;
        RECT  4.735 1.980 5.595 2.100 ;
        RECT  5.180 1.070 5.495 1.330 ;
        RECT  5.060 0.900 5.180 1.620 ;
        RECT  5.010 0.380 5.130 0.540 ;
        RECT  5.040 0.900 5.060 1.020 ;
        RECT  4.570 1.500 5.060 1.620 ;
        RECT  4.920 0.670 5.040 1.020 ;
        RECT  4.735 0.380 5.010 0.500 ;
        RECT  4.690 1.210 4.940 1.330 ;
        RECT  4.860 0.670 4.920 0.790 ;
        RECT  4.340 0.620 4.860 0.790 ;
        RECT  4.475 0.350 4.735 0.500 ;
        RECT  4.475 1.980 4.735 2.170 ;
        RECT  4.560 1.060 4.690 1.330 ;
        RECT  3.970 1.060 4.560 1.190 ;
        RECT  4.230 0.380 4.475 0.500 ;
        RECT  4.015 1.980 4.475 2.100 ;
        RECT  4.150 1.310 4.270 1.860 ;
        RECT  4.110 0.380 4.230 0.550 ;
        RECT  3.495 0.430 4.110 0.550 ;
        RECT  3.900 1.980 4.015 2.140 ;
        RECT  3.850 0.685 3.970 1.615 ;
        RECT  2.975 2.020 3.900 2.140 ;
        RECT  3.280 0.685 3.850 0.805 ;
        RECT  3.810 1.495 3.850 1.615 ;
        RECT  3.690 1.495 3.810 1.900 ;
        RECT  3.195 1.110 3.730 1.230 ;
        RECT  3.270 1.780 3.690 1.900 ;
        RECT  3.380 0.380 3.495 0.550 ;
        RECT  2.410 0.380 3.380 0.500 ;
        RECT  3.165 0.630 3.280 0.805 ;
        RECT  3.075 1.020 3.195 1.670 ;
        RECT  2.950 0.630 3.165 0.750 ;
        RECT  3.050 1.020 3.075 1.140 ;
        RECT  2.025 1.550 3.075 1.670 ;
        RECT  2.930 0.880 3.050 1.140 ;
        RECT  2.855 1.790 2.975 2.140 ;
        RECT  2.810 1.310 2.955 1.430 ;
        RECT  1.730 1.790 2.855 1.910 ;
        RECT  2.690 0.630 2.810 1.430 ;
        RECT  2.530 0.630 2.690 0.750 ;
        RECT  2.290 0.380 2.410 0.620 ;
        RECT  1.570 0.500 2.290 0.620 ;
        RECT  2.025 0.740 2.055 0.860 ;
        RECT  1.905 0.740 2.025 1.670 ;
        RECT  1.795 0.740 1.905 0.860 ;
        RECT  1.660 1.395 1.780 1.670 ;
        RECT  1.470 1.790 1.730 2.190 ;
        RECT  1.570 1.395 1.660 1.515 ;
        RECT  1.450 0.500 1.570 1.515 ;
        RECT  1.350 1.725 1.470 1.910 ;
        RECT  1.410 0.500 1.450 0.930 ;
        RECT  0.615 1.725 1.350 1.845 ;
        RECT  0.860 1.435 0.885 1.605 ;
        RECT  0.740 0.660 0.860 1.605 ;
        RECT  0.650 1.000 0.740 1.260 ;
        RECT  0.715 1.435 0.740 1.605 ;
        RECT  0.520 1.725 0.615 1.965 ;
        RECT  0.400 0.660 0.520 1.965 ;
    END
END SDFFNHX1AD
MACRO SDFFNHX2AD
    CLASS CORE ;
    FOREIGN SDFFNHX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.320 1.350 3.570 1.655 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.850 2.030 2.215 2.190 ;
        END
        AntennaGateArea 0.096 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.210 1.740 7.430 1.860 ;
        RECT  7.210 0.690 7.360 0.950 ;
        RECT  7.070 0.690 7.210 1.860 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.315 0.735 8.330 1.625 ;
        RECT  8.190 0.400 8.315 2.145 ;
        RECT  8.145 0.400 8.190 0.830 ;
        RECT  8.145 1.455 8.190 2.145 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.450 0.980 2.570 1.240 ;
        RECT  2.305 0.860 2.450 1.350 ;
        END
        AntennaGateArea 0.084 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.125 1.330 1.375 ;
        RECT  1.020 1.025 1.190 1.375 ;
        END
        AntennaGateArea 0.127 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.955 -0.210 8.400 0.210 ;
        RECT  7.785 -0.210 7.955 0.555 ;
        RECT  7.050 -0.210 7.785 0.210 ;
        RECT  6.790 -0.210 7.050 0.300 ;
        RECT  5.600 -0.210 6.790 0.210 ;
        RECT  5.340 -0.210 5.600 0.290 ;
        RECT  3.835 -0.210 5.340 0.210 ;
        RECT  3.665 -0.210 3.835 0.415 ;
        RECT  2.170 -0.210 3.665 0.210 ;
        RECT  1.910 -0.210 2.170 0.380 ;
        RECT  1.265 -0.210 1.910 0.210 ;
        RECT  1.095 -0.210 1.265 0.375 ;
        RECT  0.335 -0.210 1.095 0.210 ;
        RECT  0.165 -0.210 0.335 0.400 ;
        RECT  0.000 -0.210 0.165 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.960 2.310 8.400 2.730 ;
        RECT  7.790 1.885 7.960 2.730 ;
        RECT  7.000 2.310 7.790 2.730 ;
        RECT  6.740 2.220 7.000 2.730 ;
        RECT  5.555 2.310 6.740 2.730 ;
        RECT  5.295 2.230 5.555 2.730 ;
        RECT  4.360 2.310 5.295 2.730 ;
        RECT  4.100 2.230 4.360 2.730 ;
        RECT  2.510 2.310 4.100 2.730 ;
        RECT  2.340 2.070 2.510 2.730 ;
        RECT  1.220 2.310 2.340 2.730 ;
        RECT  0.960 1.965 1.220 2.730 ;
        RECT  0.255 2.310 0.960 2.730 ;
        RECT  0.085 1.540 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.400 2.520 ;
        LAYER M1 ;
        RECT  7.880 1.045 8.000 1.760 ;
        RECT  7.795 1.045 7.880 1.215 ;
        RECT  7.670 1.640 7.880 1.760 ;
        RECT  7.600 1.400 7.690 1.520 ;
        RECT  7.550 1.640 7.670 2.100 ;
        RECT  7.480 0.385 7.600 1.520 ;
        RECT  6.745 1.980 7.550 2.100 ;
        RECT  7.425 0.385 7.480 0.555 ;
        RECT  7.430 1.400 7.480 1.520 ;
        RECT  6.850 0.435 7.425 0.555 ;
        RECT  6.730 0.435 6.850 1.520 ;
        RECT  6.625 1.670 6.745 2.100 ;
        RECT  6.105 1.670 6.625 1.790 ;
        RECT  6.465 0.330 6.585 1.510 ;
        RECT  6.225 1.980 6.485 2.190 ;
        RECT  6.325 0.330 6.465 0.500 ;
        RECT  6.280 1.390 6.465 1.510 ;
        RECT  6.295 0.645 6.345 0.815 ;
        RECT  5.855 0.380 6.325 0.500 ;
        RECT  6.175 0.645 6.295 1.080 ;
        RECT  4.735 1.980 6.225 2.100 ;
        RECT  6.105 0.960 6.175 1.080 ;
        RECT  5.985 0.960 6.105 1.790 ;
        RECT  5.865 0.650 6.030 0.770 ;
        RECT  5.745 0.650 5.865 1.860 ;
        RECT  5.735 0.380 5.855 0.530 ;
        RECT  5.160 0.650 5.745 0.770 ;
        RECT  4.210 1.740 5.745 1.860 ;
        RECT  5.130 0.410 5.735 0.530 ;
        RECT  5.180 1.070 5.625 1.330 ;
        RECT  5.060 0.890 5.180 1.620 ;
        RECT  5.010 0.380 5.130 0.530 ;
        RECT  5.040 0.890 5.060 1.010 ;
        RECT  4.570 1.500 5.060 1.620 ;
        RECT  4.920 0.650 5.040 1.010 ;
        RECT  4.735 0.380 5.010 0.500 ;
        RECT  4.690 1.190 4.940 1.310 ;
        RECT  4.860 0.650 4.920 0.770 ;
        RECT  4.340 0.620 4.860 0.770 ;
        RECT  4.475 0.350 4.735 0.500 ;
        RECT  4.475 1.980 4.735 2.190 ;
        RECT  4.560 1.060 4.690 1.310 ;
        RECT  3.970 1.060 4.560 1.190 ;
        RECT  4.150 0.380 4.475 0.500 ;
        RECT  4.015 1.980 4.475 2.100 ;
        RECT  4.090 1.340 4.210 1.860 ;
        RECT  4.030 0.380 4.150 0.655 ;
        RECT  3.545 0.535 4.030 0.655 ;
        RECT  3.900 1.980 4.015 2.140 ;
        RECT  3.850 0.775 3.970 1.470 ;
        RECT  2.865 2.020 3.900 2.140 ;
        RECT  3.305 0.775 3.850 0.895 ;
        RECT  3.810 1.350 3.850 1.470 ;
        RECT  3.690 1.350 3.810 1.900 ;
        RECT  3.195 1.110 3.730 1.230 ;
        RECT  3.080 1.780 3.690 1.900 ;
        RECT  3.425 0.380 3.545 0.655 ;
        RECT  2.410 0.380 3.425 0.500 ;
        RECT  3.185 0.630 3.305 0.895 ;
        RECT  3.075 1.060 3.195 1.660 ;
        RECT  2.950 0.630 3.185 0.750 ;
        RECT  3.050 1.060 3.075 1.180 ;
        RECT  2.145 1.540 3.075 1.660 ;
        RECT  2.930 0.920 3.050 1.180 ;
        RECT  2.810 1.300 2.955 1.420 ;
        RECT  2.745 1.790 2.865 2.140 ;
        RECT  2.690 0.630 2.810 1.420 ;
        RECT  1.730 1.790 2.745 1.910 ;
        RECT  2.530 0.630 2.690 0.750 ;
        RECT  2.290 0.380 2.410 0.620 ;
        RECT  1.570 0.500 2.290 0.620 ;
        RECT  2.055 1.425 2.145 1.660 ;
        RECT  1.935 0.740 2.055 1.660 ;
        RECT  1.795 0.740 1.935 0.860 ;
        RECT  1.660 1.395 1.780 1.670 ;
        RECT  1.470 1.790 1.730 2.190 ;
        RECT  1.570 1.395 1.660 1.515 ;
        RECT  1.450 0.500 1.570 1.515 ;
        RECT  1.350 1.725 1.470 1.910 ;
        RECT  1.410 0.500 1.450 0.930 ;
        RECT  0.615 1.725 1.350 1.845 ;
        RECT  0.860 1.435 0.885 1.605 ;
        RECT  0.715 0.660 0.860 1.605 ;
        RECT  0.650 1.000 0.715 1.260 ;
        RECT  0.520 1.725 0.615 2.065 ;
        RECT  0.400 0.660 0.520 2.065 ;
    END
END SDFFNHX2AD
MACRO SDFFNHX4AD
    CLASS CORE ;
    FOREIGN SDFFNHX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.125 1.410 4.505 1.610 ;
        END
        AntennaGateArea 0.076 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.525 2.020 3.785 2.190 ;
        RECT  2.805 2.020 3.525 2.140 ;
        RECT  2.525 2.020 2.805 2.190 ;
        END
        AntennaGateArea 0.124 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.715 1.750 9.945 1.900 ;
        RECT  9.715 0.735 9.800 0.905 ;
        RECT  9.585 0.735 9.715 1.900 ;
        RECT  9.405 1.750 9.585 1.900 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.790 1.005 10.850 1.515 ;
        RECT  10.660 0.410 10.790 2.090 ;
        RECT  10.585 0.410 10.660 0.840 ;
        RECT  10.585 1.400 10.660 2.090 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.820 0.865 3.030 1.390 ;
        END
        AntennaGateArea 0.138 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.315 1.100 1.610 1.375 ;
        END
        AntennaGateArea 0.167 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.115 -0.210 11.200 0.210 ;
        RECT  10.945 -0.210 11.115 0.810 ;
        RECT  10.370 -0.210 10.945 0.210 ;
        RECT  10.250 -0.210 10.370 0.805 ;
        RECT  9.455 -0.210 10.250 0.210 ;
        RECT  9.195 -0.210 9.455 0.300 ;
        RECT  8.650 -0.210 9.195 0.210 ;
        RECT  8.390 -0.210 8.650 0.240 ;
        RECT  6.980 -0.210 8.390 0.210 ;
        RECT  6.720 -0.210 6.980 0.260 ;
        RECT  4.950 -0.210 6.720 0.210 ;
        RECT  4.430 -0.210 4.950 0.260 ;
        RECT  2.670 -0.210 4.430 0.210 ;
        RECT  2.550 -0.210 2.670 0.500 ;
        RECT  1.515 -0.210 2.550 0.210 ;
        RECT  1.345 -0.210 1.515 0.885 ;
        RECT  0.285 -0.210 1.345 0.210 ;
        RECT  0.165 -0.210 0.285 0.920 ;
        RECT  0.000 -0.210 0.165 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.090 2.310 11.200 2.730 ;
        RECT  10.970 1.505 11.090 2.730 ;
        RECT  10.325 2.310 10.970 2.730 ;
        RECT  10.155 2.265 10.325 2.730 ;
        RECT  9.520 2.310 10.155 2.730 ;
        RECT  9.350 2.265 9.520 2.730 ;
        RECT  8.770 2.310 9.350 2.730 ;
        RECT  8.510 2.220 8.770 2.730 ;
        RECT  7.130 2.310 8.510 2.730 ;
        RECT  6.960 2.265 7.130 2.730 ;
        RECT  6.185 2.310 6.960 2.730 ;
        RECT  5.925 2.290 6.185 2.730 ;
        RECT  5.040 2.310 5.925 2.730 ;
        RECT  4.780 2.260 5.040 2.730 ;
        RECT  3.165 2.310 4.780 2.730 ;
        RECT  2.905 2.260 3.165 2.730 ;
        RECT  1.585 2.310 2.905 2.730 ;
        RECT  1.325 2.190 1.585 2.730 ;
        RECT  0.615 2.310 1.325 2.730 ;
        RECT  0.445 1.630 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.200 2.520 ;
        LAYER M1 ;
        RECT  10.280 0.990 10.540 1.250 ;
        RECT  10.160 0.990 10.280 2.140 ;
        RECT  9.090 2.020 10.160 2.140 ;
        RECT  9.920 0.420 10.040 1.545 ;
        RECT  9.440 0.420 9.920 0.540 ;
        RECT  9.835 1.375 9.920 1.545 ;
        RECT  9.320 0.420 9.440 1.575 ;
        RECT  8.970 1.750 9.090 2.140 ;
        RECT  8.965 0.380 9.085 1.620 ;
        RECT  8.845 1.750 8.970 1.900 ;
        RECT  7.700 0.380 8.965 0.500 ;
        RECT  8.725 0.690 8.845 1.900 ;
        RECT  7.945 1.480 8.725 1.600 ;
        RECT  8.135 1.780 8.305 1.950 ;
        RECT  7.500 0.620 8.270 0.740 ;
        RECT  7.620 1.780 8.135 1.900 ;
        RECT  7.880 1.480 7.945 1.650 ;
        RECT  7.740 0.865 7.880 1.650 ;
        RECT  7.540 2.020 7.800 2.190 ;
        RECT  7.620 0.865 7.740 0.985 ;
        RECT  7.440 0.330 7.700 0.500 ;
        RECT  7.500 1.690 7.620 1.900 ;
        RECT  5.435 2.020 7.540 2.140 ;
        RECT  7.380 0.620 7.500 1.900 ;
        RECT  6.395 0.380 7.440 0.500 ;
        RECT  7.200 0.620 7.380 0.790 ;
        RECT  7.090 1.780 7.380 1.900 ;
        RECT  6.850 0.950 7.245 1.070 ;
        RECT  6.970 1.215 7.090 1.900 ;
        RECT  5.060 1.780 6.970 1.900 ;
        RECT  6.730 0.900 6.850 1.660 ;
        RECT  6.435 0.900 6.730 1.020 ;
        RECT  5.370 1.540 6.730 1.660 ;
        RECT  6.475 1.160 6.595 1.420 ;
        RECT  5.765 1.300 6.475 1.420 ;
        RECT  6.315 0.640 6.435 1.020 ;
        RECT  5.875 0.360 6.395 0.500 ;
        RECT  5.640 0.640 6.315 0.760 ;
        RECT  2.910 0.380 5.875 0.500 ;
        RECT  5.305 1.265 5.765 1.420 ;
        RECT  5.175 2.020 5.435 2.190 ;
        RECT  5.185 0.620 5.305 1.420 ;
        RECT  4.820 0.620 5.185 0.740 ;
        RECT  4.030 2.020 5.175 2.140 ;
        RECT  4.940 1.150 5.060 1.900 ;
        RECT  4.700 0.620 4.820 1.900 ;
        RECT  3.650 0.620 4.700 0.740 ;
        RECT  4.150 1.780 4.700 1.900 ;
        RECT  4.460 0.965 4.580 1.280 ;
        RECT  4.005 0.965 4.460 1.085 ;
        RECT  3.910 1.780 4.030 2.140 ;
        RECT  3.885 0.965 4.005 1.650 ;
        RECT  2.405 1.780 3.910 1.900 ;
        RECT  3.410 0.965 3.885 1.085 ;
        RECT  2.550 1.525 3.885 1.650 ;
        RECT  3.290 1.265 3.765 1.385 ;
        RECT  3.170 0.620 3.290 1.385 ;
        RECT  3.030 0.620 3.170 0.740 ;
        RECT  2.790 0.380 2.910 0.740 ;
        RECT  2.430 0.620 2.790 0.740 ;
        RECT  2.335 1.290 2.550 1.650 ;
        RECT  2.310 0.385 2.430 0.740 ;
        RECT  2.285 1.780 2.405 2.140 ;
        RECT  2.190 1.290 2.335 1.410 ;
        RECT  1.850 0.385 2.310 0.505 ;
        RECT  1.845 2.020 2.285 2.140 ;
        RECT  2.070 0.675 2.190 1.410 ;
        RECT  2.025 1.550 2.145 1.810 ;
        RECT  1.850 1.550 2.025 1.670 ;
        RECT  1.730 0.385 1.850 1.670 ;
        RECT  1.725 1.930 1.845 2.140 ;
        RECT  0.975 1.930 1.725 2.050 ;
        RECT  1.155 1.515 1.250 1.685 ;
        RECT  1.035 0.680 1.155 1.685 ;
        RECT  0.985 0.680 1.035 1.190 ;
        RECT  0.770 1.055 0.985 1.190 ;
        RECT  0.910 1.880 0.975 2.050 ;
        RECT  0.780 1.390 0.910 2.050 ;
        RECT  0.530 1.390 0.780 1.510 ;
        RECT  0.650 1.000 0.770 1.260 ;
        RECT  0.530 0.415 0.670 0.845 ;
        RECT  0.500 0.415 0.530 1.510 ;
        RECT  0.405 0.640 0.500 1.510 ;
        RECT  0.255 1.390 0.405 1.510 ;
        RECT  0.085 1.390 0.255 1.975 ;
    END
END SDFFNHX4AD
MACRO SDFFNHX8AD
    CLASS CORE ;
    FOREIGN SDFFNHX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.960 1.265 5.340 1.610 ;
        END
        AntennaGateArea 0.113 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.870 0.770 3.030 1.150 ;
        RECT  2.770 1.030 2.870 1.150 ;
        END
        AntennaGateArea 0.165 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.995 0.660 13.090 0.830 ;
        RECT  12.995 1.780 13.080 1.900 ;
        RECT  12.865 0.660 12.995 1.900 ;
        RECT  12.820 1.330 12.865 1.900 ;
        RECT  12.485 1.330 12.820 1.780 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.675 1.000 14.910 1.625 ;
        RECT  14.505 0.380 14.675 2.145 ;
        RECT  14.425 0.665 14.505 1.625 ;
        RECT  13.955 0.665 14.425 0.915 ;
        RECT  13.955 1.375 14.425 1.625 ;
        RECT  13.785 0.410 13.955 0.915 ;
        RECT  13.785 1.375 13.955 2.155 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.455 1.095 3.885 1.265 ;
        RECT  3.150 1.095 3.455 1.375 ;
        END
        AntennaGateArea 0.262 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.080 2.065 1.260 ;
        RECT  1.750 1.080 1.890 1.655 ;
        END
        AntennaGateArea 0.275 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.035 -0.210 15.120 0.210 ;
        RECT  14.865 -0.210 15.035 0.810 ;
        RECT  14.315 -0.210 14.865 0.210 ;
        RECT  14.145 -0.210 14.315 0.490 ;
        RECT  13.570 -0.210 14.145 0.210 ;
        RECT  13.450 -0.210 13.570 0.805 ;
        RECT  12.755 -0.210 13.450 0.210 ;
        RECT  12.495 -0.210 12.755 0.260 ;
        RECT  9.820 -0.210 12.495 0.210 ;
        RECT  9.650 -0.210 9.820 0.260 ;
        RECT  9.060 -0.210 9.650 0.210 ;
        RECT  8.890 -0.210 9.060 0.260 ;
        RECT  8.260 -0.210 8.890 0.210 ;
        RECT  8.000 -0.210 8.260 0.260 ;
        RECT  6.095 -0.210 8.000 0.210 ;
        RECT  5.575 -0.210 6.095 0.260 ;
        RECT  3.860 -0.210 5.575 0.210 ;
        RECT  3.600 -0.210 3.860 0.380 ;
        RECT  3.095 -0.210 3.600 0.210 ;
        RECT  2.835 -0.210 3.095 0.380 ;
        RECT  1.970 -0.210 2.835 0.210 ;
        RECT  1.800 -0.210 1.970 0.825 ;
        RECT  1.030 -0.210 1.800 0.210 ;
        RECT  0.860 -0.210 1.030 0.845 ;
        RECT  0.310 -0.210 0.860 0.210 ;
        RECT  0.140 -0.210 0.310 0.845 ;
        RECT  0.000 -0.210 0.140 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.035 2.310 15.120 2.730 ;
        RECT  14.865 1.775 15.035 2.730 ;
        RECT  14.315 2.310 14.865 2.730 ;
        RECT  14.145 1.765 14.315 2.730 ;
        RECT  13.525 2.310 14.145 2.730 ;
        RECT  13.355 2.265 13.525 2.730 ;
        RECT  12.655 2.310 13.355 2.730 ;
        RECT  12.485 2.265 12.655 2.730 ;
        RECT  9.545 2.310 12.485 2.730 ;
        RECT  9.285 2.005 9.545 2.730 ;
        RECT  8.805 2.310 9.285 2.730 ;
        RECT  8.545 2.265 8.805 2.730 ;
        RECT  7.260 2.310 8.545 2.730 ;
        RECT  7.000 2.290 7.260 2.730 ;
        RECT  5.925 2.310 7.000 2.730 ;
        RECT  5.665 2.260 5.925 2.730 ;
        RECT  4.220 2.310 5.665 2.730 ;
        RECT  3.960 2.140 4.220 2.730 ;
        RECT  3.460 2.310 3.960 2.730 ;
        RECT  3.200 2.140 3.460 2.730 ;
        RECT  2.040 2.310 3.200 2.730 ;
        RECT  1.780 2.190 2.040 2.730 ;
        RECT  0.975 2.310 1.780 2.730 ;
        RECT  0.805 1.630 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.630 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 15.120 2.520 ;
        LAYER M1 ;
        RECT  13.585 1.090 14.245 1.210 ;
        RECT  13.465 1.090 13.585 2.140 ;
        RECT  12.100 2.020 13.465 2.140 ;
        RECT  13.210 0.345 13.330 1.590 ;
        RECT  12.980 0.345 13.210 0.540 ;
        RECT  13.140 1.330 13.210 1.590 ;
        RECT  12.640 0.420 12.980 0.540 ;
        RECT  12.520 0.420 12.640 1.155 ;
        RECT  12.280 0.380 12.400 1.225 ;
        RECT  7.435 0.380 12.280 0.500 ;
        RECT  12.165 1.105 12.280 1.225 ;
        RECT  12.045 1.105 12.165 1.555 ;
        RECT  11.990 0.660 12.160 0.985 ;
        RECT  11.925 1.755 12.100 2.140 ;
        RECT  11.925 0.865 11.990 0.985 ;
        RECT  11.805 0.865 11.925 2.140 ;
        RECT  9.835 0.620 11.865 0.740 ;
        RECT  10.440 0.865 11.805 0.985 ;
        RECT  11.395 2.020 11.805 2.140 ;
        RECT  11.565 1.505 11.685 1.765 ;
        RECT  9.835 1.505 11.565 1.625 ;
        RECT  11.135 1.745 11.395 2.140 ;
        RECT  10.670 1.745 11.135 1.865 ;
        RECT  10.410 1.745 10.670 2.125 ;
        RECT  9.860 1.755 10.120 2.190 ;
        RECT  8.640 1.755 9.860 1.875 ;
        RECT  9.715 0.620 9.835 1.625 ;
        RECT  8.465 0.620 9.715 0.740 ;
        RECT  8.335 1.505 9.715 1.625 ;
        RECT  7.965 1.025 9.340 1.195 ;
        RECT  8.520 1.755 8.640 2.140 ;
        RECT  6.435 2.020 8.520 2.140 ;
        RECT  8.165 1.505 8.335 1.900 ;
        RECT  6.095 1.780 8.165 1.900 ;
        RECT  7.845 0.900 7.965 1.660 ;
        RECT  7.395 0.900 7.845 1.020 ;
        RECT  6.370 1.540 7.845 1.660 ;
        RECT  7.590 1.160 7.710 1.420 ;
        RECT  6.730 1.300 7.590 1.420 ;
        RECT  6.915 0.360 7.435 0.500 ;
        RECT  7.235 0.640 7.395 1.020 ;
        RECT  6.675 0.640 7.235 0.760 ;
        RECT  4.355 0.380 6.915 0.500 ;
        RECT  6.340 1.210 6.730 1.420 ;
        RECT  6.175 2.020 6.435 2.190 ;
        RECT  6.220 0.620 6.340 1.420 ;
        RECT  5.855 0.620 6.220 0.740 ;
        RECT  4.865 2.020 6.175 2.140 ;
        RECT  5.975 1.150 6.095 1.900 ;
        RECT  5.735 0.620 5.855 1.900 ;
        RECT  4.485 0.620 5.735 0.740 ;
        RECT  4.985 1.780 5.735 1.900 ;
        RECT  4.840 0.965 5.615 1.085 ;
        RECT  4.745 1.900 4.865 2.140 ;
        RECT  4.720 0.965 4.840 1.780 ;
        RECT  2.860 1.900 4.745 2.020 ;
        RECT  4.690 0.965 4.720 1.085 ;
        RECT  3.050 1.655 4.720 1.780 ;
        RECT  4.430 0.930 4.690 1.085 ;
        RECT  4.125 1.415 4.600 1.535 ;
        RECT  4.235 0.380 4.355 0.620 ;
        RECT  4.125 0.740 4.240 0.860 ;
        RECT  2.305 0.500 4.235 0.620 ;
        RECT  4.005 0.740 4.125 1.535 ;
        RECT  3.220 0.740 4.005 0.860 ;
        RECT  3.580 1.415 4.005 1.535 ;
        RECT  3.005 1.610 3.050 1.780 ;
        RECT  2.790 1.290 3.005 1.780 ;
        RECT  2.740 1.900 2.860 2.140 ;
        RECT  2.645 1.290 2.790 1.410 ;
        RECT  2.300 2.020 2.740 2.140 ;
        RECT  2.645 0.745 2.715 0.865 ;
        RECT  2.525 0.745 2.645 1.410 ;
        RECT  2.480 1.550 2.600 1.810 ;
        RECT  2.455 0.745 2.525 0.865 ;
        RECT  2.305 1.550 2.480 1.670 ;
        RECT  2.185 0.500 2.305 1.670 ;
        RECT  2.180 1.930 2.300 2.140 ;
        RECT  1.335 1.930 2.180 2.050 ;
        RECT  1.445 0.380 1.615 1.685 ;
        RECT  1.440 0.380 1.445 1.190 ;
        RECT  1.155 1.055 1.440 1.190 ;
        RECT  1.270 1.880 1.335 2.050 ;
        RECT  1.140 1.390 1.270 2.050 ;
        RECT  0.775 1.000 1.155 1.260 ;
        RECT  0.655 1.390 1.140 1.510 ;
        RECT  0.615 0.385 0.655 1.510 ;
        RECT  0.525 0.385 0.615 1.975 ;
        RECT  0.445 1.390 0.525 1.975 ;
    END
END SDFFNHX8AD
MACRO SDFFNSRHX1AD
    CLASS CORE ;
    FOREIGN SDFFNSRHX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.725 1.080 4.985 1.375 ;
        END
        AntennaGateArea 0.115 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.795 0.860 3.010 1.120 ;
        RECT  2.545 0.860 2.795 1.030 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.145 0.865 3.315 1.420 ;
        RECT  2.660 1.300 3.145 1.420 ;
        RECT  2.540 1.160 2.660 1.420 ;
        END
        AntennaGateArea 0.096 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.185 1.020 9.305 1.280 ;
        RECT  7.815 1.080 9.185 1.200 ;
        RECT  7.585 1.080 7.815 1.330 ;
        END
        AntennaGateArea 0.108 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.470 1.425 10.595 1.710 ;
        RECT  10.350 0.910 10.470 1.710 ;
        RECT  10.130 0.910 10.350 1.030 ;
        END
        AntennaDiffArea 0.192 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.650 1.145 11.690 1.375 ;
        RECT  11.530 0.645 11.650 1.915 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.920 1.895 1.375 ;
        END
        AntennaGateArea 0.061 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.955 0.490 1.375 ;
        END
        AntennaGateArea 0.118 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.340 -0.210 11.760 0.210 ;
        RECT  11.080 -0.210 11.340 0.310 ;
        RECT  10.690 -0.210 11.080 0.210 ;
        RECT  10.430 -0.210 10.690 0.310 ;
        RECT  9.950 -0.210 10.430 0.210 ;
        RECT  9.690 -0.210 9.950 0.310 ;
        RECT  8.045 -0.210 9.690 0.210 ;
        RECT  7.785 -0.210 8.045 0.310 ;
        RECT  6.740 -0.210 7.785 0.210 ;
        RECT  6.480 -0.210 6.740 0.310 ;
        RECT  4.950 -0.210 6.480 0.210 ;
        RECT  4.520 -0.210 4.950 0.255 ;
        RECT  3.720 -0.210 4.520 0.210 ;
        RECT  3.290 -0.210 3.720 0.255 ;
        RECT  1.655 -0.210 3.290 0.210 ;
        RECT  1.395 -0.210 1.655 0.310 ;
        RECT  0.545 -0.210 1.395 0.210 ;
        RECT  0.425 -0.210 0.545 0.380 ;
        RECT  0.000 -0.210 0.425 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.275 2.310 11.760 2.730 ;
        RECT  10.845 2.150 11.275 2.730 ;
        RECT  9.490 2.310 10.845 2.730 ;
        RECT  9.230 2.230 9.490 2.730 ;
        RECT  7.830 2.310 9.230 2.730 ;
        RECT  7.660 2.265 7.830 2.730 ;
        RECT  7.245 2.310 7.660 2.730 ;
        RECT  6.985 2.220 7.245 2.730 ;
        RECT  6.305 2.310 6.985 2.730 ;
        RECT  6.045 2.220 6.305 2.730 ;
        RECT  4.800 2.310 6.045 2.730 ;
        RECT  4.280 2.220 4.800 2.730 ;
        RECT  3.670 2.310 4.280 2.730 ;
        RECT  3.410 2.260 3.670 2.730 ;
        RECT  1.885 2.310 3.410 2.730 ;
        RECT  1.625 2.210 1.885 2.730 ;
        RECT  0.560 2.310 1.625 2.730 ;
        RECT  0.390 1.925 0.560 2.730 ;
        RECT  0.000 2.310 0.390 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.760 2.520 ;
        LAYER M1 ;
        RECT  11.245 1.065 11.410 1.235 ;
        RECT  11.125 0.430 11.245 2.030 ;
        RECT  10.330 0.430 11.125 0.550 ;
        RECT  10.980 1.065 11.125 1.235 ;
        RECT  10.390 1.910 11.125 2.030 ;
        RECT  10.835 0.670 11.005 0.905 ;
        RECT  10.835 1.410 11.005 1.580 ;
        RECT  10.715 0.670 10.835 1.580 ;
        RECT  10.590 0.670 10.715 1.260 ;
        RECT  9.790 0.670 10.590 0.790 ;
        RECT  10.130 1.910 10.390 2.045 ;
        RECT  10.070 0.380 10.330 0.550 ;
        RECT  10.110 1.150 10.230 1.780 ;
        RECT  8.635 1.925 10.130 2.045 ;
        RECT  9.550 1.150 10.110 1.270 ;
        RECT  9.005 0.430 10.070 0.550 ;
        RECT  9.710 1.390 9.970 1.580 ;
        RECT  9.670 0.670 9.790 0.960 ;
        RECT  8.915 1.460 9.710 1.580 ;
        RECT  9.430 0.780 9.550 1.270 ;
        RECT  8.715 0.780 9.430 0.900 ;
        RECT  8.835 0.355 9.005 0.550 ;
        RECT  8.795 1.460 8.915 1.800 ;
        RECT  8.345 1.680 8.795 1.800 ;
        RECT  8.595 0.430 8.715 0.900 ;
        RECT  8.425 0.430 8.595 0.550 ;
        RECT  8.085 1.440 8.515 1.560 ;
        RECT  8.255 2.020 8.515 2.180 ;
        RECT  7.310 0.705 8.475 0.875 ;
        RECT  8.165 0.340 8.425 0.550 ;
        RECT  8.225 1.680 8.345 1.870 ;
        RECT  7.675 2.020 8.255 2.140 ;
        RECT  7.775 1.730 8.225 1.870 ;
        RECT  6.120 0.430 8.165 0.550 ;
        RECT  7.965 1.440 8.085 1.610 ;
        RECT  7.310 1.490 7.965 1.610 ;
        RECT  6.755 1.730 7.775 1.850 ;
        RECT  7.555 1.980 7.675 2.140 ;
        RECT  6.725 1.980 7.555 2.100 ;
        RECT  7.190 0.705 7.310 1.610 ;
        RECT  6.875 1.395 7.190 1.515 ;
        RECT  6.975 0.675 7.055 0.795 ;
        RECT  6.855 0.675 6.975 1.275 ;
        RECT  4.555 0.675 6.855 0.795 ;
        RECT  6.755 1.155 6.855 1.275 ;
        RECT  6.635 1.155 6.755 1.850 ;
        RECT  6.465 1.980 6.725 2.185 ;
        RECT  6.515 0.915 6.705 1.035 ;
        RECT  6.395 0.915 6.515 1.850 ;
        RECT  5.365 1.980 6.465 2.100 ;
        RECT  5.675 0.915 6.395 1.035 ;
        RECT  5.605 1.550 6.395 1.670 ;
        RECT  5.860 0.330 6.120 0.550 ;
        RECT  4.605 0.430 5.860 0.550 ;
        RECT  5.485 1.550 5.605 1.810 ;
        RECT  5.365 1.000 5.395 1.260 ;
        RECT  5.245 1.000 5.365 2.100 ;
        RECT  4.160 1.980 5.245 2.100 ;
        RECT  4.160 1.740 5.125 1.860 ;
        RECT  4.485 0.380 4.605 0.550 ;
        RECT  4.435 0.675 4.555 1.620 ;
        RECT  1.895 0.380 4.485 0.500 ;
        RECT  4.280 1.500 4.435 1.620 ;
        RECT  4.195 0.620 4.315 1.230 ;
        RECT  3.570 0.620 4.195 0.740 ;
        RECT  4.160 1.105 4.195 1.230 ;
        RECT  4.040 1.105 4.160 1.860 ;
        RECT  4.040 1.980 4.160 2.140 ;
        RECT  3.920 0.860 4.075 0.980 ;
        RECT  2.135 2.020 4.040 2.140 ;
        RECT  3.800 0.860 3.920 1.900 ;
        RECT  2.375 1.780 3.800 1.900 ;
        RECT  3.450 0.620 3.570 1.660 ;
        RECT  2.605 0.620 3.450 0.740 ;
        RECT  2.590 1.540 3.450 1.660 ;
        RECT  2.375 0.860 2.425 1.120 ;
        RECT  2.135 0.620 2.420 0.740 ;
        RECT  2.255 0.860 2.375 1.900 ;
        RECT  2.015 0.620 2.135 1.745 ;
        RECT  2.015 1.960 2.135 2.140 ;
        RECT  1.435 1.960 2.015 2.080 ;
        RECT  1.775 0.380 1.895 0.740 ;
        RECT  1.025 0.620 1.775 0.740 ;
        RECT  1.435 0.860 1.505 0.980 ;
        RECT  1.315 0.860 1.435 2.080 ;
        RECT  1.245 0.860 1.315 1.385 ;
        RECT  0.785 0.380 1.275 0.500 ;
        RECT  1.155 1.125 1.245 1.385 ;
        RECT  1.025 1.770 1.165 2.030 ;
        RECT  0.905 0.620 1.025 2.030 ;
        RECT  0.665 0.380 0.785 0.835 ;
        RECT  0.270 0.715 0.665 0.835 ;
        RECT  0.220 0.665 0.270 0.835 ;
        RECT  0.220 1.495 0.270 1.665 ;
        RECT  0.100 0.665 0.220 1.665 ;
    END
END SDFFNSRHX1AD
MACRO SDFFNSRHX2AD
    CLASS CORE ;
    FOREIGN SDFFNSRHX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.675 1.010 5.070 1.375 ;
        END
        AntennaGateArea 0.137 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.795 0.860 3.010 1.120 ;
        RECT  2.545 0.860 2.795 1.030 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.145 0.865 3.315 1.420 ;
        RECT  2.660 1.300 3.145 1.420 ;
        RECT  2.540 1.160 2.660 1.420 ;
        END
        AntennaGateArea 0.096 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.165 1.020 9.285 1.280 ;
        RECT  7.815 1.080 9.165 1.200 ;
        RECT  7.585 1.080 7.815 1.330 ;
        END
        AntennaGateArea 0.138 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.470 1.425 10.595 1.710 ;
        RECT  10.350 0.910 10.470 1.710 ;
        RECT  10.130 0.910 10.350 1.030 ;
        END
        AntennaDiffArea 0.192 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.530 0.330 11.690 1.915 ;
        END
        AntennaDiffArea 0.368 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.920 1.895 1.375 ;
        END
        AntennaGateArea 0.088 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.040 0.770 1.375 ;
        END
        AntennaGateArea 0.127 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.290 -0.210 11.760 0.210 ;
        RECT  11.030 -0.210 11.290 0.310 ;
        RECT  10.690 -0.210 11.030 0.210 ;
        RECT  10.430 -0.210 10.690 0.310 ;
        RECT  9.950 -0.210 10.430 0.210 ;
        RECT  9.690 -0.210 9.950 0.310 ;
        RECT  8.000 -0.210 9.690 0.210 ;
        RECT  7.830 -0.210 8.000 0.290 ;
        RECT  6.740 -0.210 7.830 0.210 ;
        RECT  6.480 -0.210 6.740 0.310 ;
        RECT  4.900 -0.210 6.480 0.210 ;
        RECT  4.470 -0.210 4.900 0.255 ;
        RECT  3.740 -0.210 4.470 0.210 ;
        RECT  3.310 -0.210 3.740 0.255 ;
        RECT  1.655 -0.210 3.310 0.210 ;
        RECT  1.395 -0.210 1.655 0.310 ;
        RECT  0.545 -0.210 1.395 0.210 ;
        RECT  0.425 -0.210 0.545 0.400 ;
        RECT  0.000 -0.210 0.425 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.255 2.310 11.760 2.730 ;
        RECT  10.825 2.165 11.255 2.730 ;
        RECT  9.445 2.310 10.825 2.730 ;
        RECT  9.275 2.265 9.445 2.730 ;
        RECT  7.800 2.310 9.275 2.730 ;
        RECT  7.630 2.265 7.800 2.730 ;
        RECT  7.080 2.310 7.630 2.730 ;
        RECT  6.910 2.265 7.080 2.730 ;
        RECT  6.305 2.310 6.910 2.730 ;
        RECT  6.045 2.220 6.305 2.730 ;
        RECT  4.800 2.310 6.045 2.730 ;
        RECT  4.280 2.220 4.800 2.730 ;
        RECT  3.670 2.310 4.280 2.730 ;
        RECT  3.410 2.260 3.670 2.730 ;
        RECT  1.935 2.310 3.410 2.730 ;
        RECT  1.675 2.240 1.935 2.730 ;
        RECT  0.560 2.310 1.675 2.730 ;
        RECT  0.390 1.975 0.560 2.730 ;
        RECT  0.000 2.310 0.390 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.760 2.520 ;
        LAYER M1 ;
        RECT  11.245 1.065 11.410 1.235 ;
        RECT  11.125 0.430 11.245 2.045 ;
        RECT  10.330 0.430 11.125 0.550 ;
        RECT  10.980 1.065 11.125 1.235 ;
        RECT  8.595 1.925 11.125 2.045 ;
        RECT  10.835 0.670 11.005 0.905 ;
        RECT  10.835 1.410 11.005 1.580 ;
        RECT  10.715 0.670 10.835 1.580 ;
        RECT  10.590 0.670 10.715 1.260 ;
        RECT  9.790 0.670 10.590 0.790 ;
        RECT  10.070 0.380 10.330 0.550 ;
        RECT  10.110 1.150 10.230 1.780 ;
        RECT  9.550 1.150 10.110 1.270 ;
        RECT  8.985 0.430 10.070 0.550 ;
        RECT  9.710 1.390 9.970 1.560 ;
        RECT  9.670 0.670 9.790 0.960 ;
        RECT  8.905 1.440 9.710 1.560 ;
        RECT  9.430 0.780 9.550 1.270 ;
        RECT  8.695 0.780 9.430 0.900 ;
        RECT  8.815 0.355 8.985 0.550 ;
        RECT  8.785 1.440 8.905 1.800 ;
        RECT  8.345 1.680 8.785 1.800 ;
        RECT  8.575 0.430 8.695 0.900 ;
        RECT  8.405 0.430 8.575 0.550 ;
        RECT  8.085 1.440 8.515 1.560 ;
        RECT  8.195 0.670 8.455 0.875 ;
        RECT  8.145 0.330 8.405 0.550 ;
        RECT  8.225 1.680 8.345 1.880 ;
        RECT  8.045 2.020 8.305 2.190 ;
        RECT  7.755 1.730 8.225 1.880 ;
        RECT  7.310 0.705 8.195 0.875 ;
        RECT  6.120 0.430 8.145 0.550 ;
        RECT  7.965 1.440 8.085 1.610 ;
        RECT  7.675 2.020 8.045 2.140 ;
        RECT  7.310 1.490 7.965 1.610 ;
        RECT  6.735 1.730 7.755 1.850 ;
        RECT  7.555 1.980 7.675 2.140 ;
        RECT  6.705 1.980 7.555 2.100 ;
        RECT  7.190 0.705 7.310 1.610 ;
        RECT  6.855 1.395 7.190 1.515 ;
        RECT  6.975 0.675 7.055 0.795 ;
        RECT  6.855 0.675 6.975 1.275 ;
        RECT  4.555 0.675 6.855 0.795 ;
        RECT  6.735 1.155 6.855 1.275 ;
        RECT  6.615 1.155 6.735 1.850 ;
        RECT  6.495 0.915 6.705 1.035 ;
        RECT  6.445 1.980 6.705 2.185 ;
        RECT  6.375 0.915 6.495 1.850 ;
        RECT  5.365 1.980 6.445 2.100 ;
        RECT  5.675 0.915 6.375 1.035 ;
        RECT  5.605 1.550 6.375 1.670 ;
        RECT  5.860 0.330 6.120 0.550 ;
        RECT  4.605 0.430 5.860 0.550 ;
        RECT  5.485 1.550 5.605 1.810 ;
        RECT  5.365 1.000 5.395 1.260 ;
        RECT  5.245 1.000 5.365 2.100 ;
        RECT  4.160 1.980 5.245 2.100 ;
        RECT  4.160 1.740 5.125 1.860 ;
        RECT  4.485 0.380 4.605 0.550 ;
        RECT  4.435 0.675 4.555 1.620 ;
        RECT  1.895 0.380 4.485 0.500 ;
        RECT  4.280 1.500 4.435 1.620 ;
        RECT  4.195 0.620 4.315 1.230 ;
        RECT  3.570 0.620 4.195 0.740 ;
        RECT  4.160 1.105 4.195 1.230 ;
        RECT  4.040 1.105 4.160 1.860 ;
        RECT  4.040 1.980 4.160 2.140 ;
        RECT  3.920 0.860 4.075 0.980 ;
        RECT  2.135 2.020 4.040 2.140 ;
        RECT  3.800 0.860 3.920 1.900 ;
        RECT  2.375 1.780 3.800 1.900 ;
        RECT  3.450 0.620 3.570 1.660 ;
        RECT  2.605 0.620 3.450 0.740 ;
        RECT  2.590 1.540 3.450 1.660 ;
        RECT  2.375 0.860 2.425 1.120 ;
        RECT  2.135 0.620 2.420 0.740 ;
        RECT  2.255 0.860 2.375 1.900 ;
        RECT  2.015 0.620 2.135 1.745 ;
        RECT  2.015 1.960 2.135 2.140 ;
        RECT  1.435 1.960 2.015 2.080 ;
        RECT  1.775 0.380 1.895 0.740 ;
        RECT  1.025 0.620 1.775 0.740 ;
        RECT  1.435 0.860 1.505 0.980 ;
        RECT  1.315 0.860 1.435 2.080 ;
        RECT  1.245 0.860 1.315 1.385 ;
        RECT  0.785 0.380 1.275 0.500 ;
        RECT  1.155 1.125 1.245 1.385 ;
        RECT  1.025 1.760 1.165 2.020 ;
        RECT  0.905 0.620 1.025 2.020 ;
        RECT  0.665 0.380 0.785 0.835 ;
        RECT  0.270 0.715 0.665 0.835 ;
        RECT  0.220 0.665 0.270 0.835 ;
        RECT  0.220 1.510 0.270 1.680 ;
        RECT  0.100 0.665 0.220 1.680 ;
    END
END SDFFNSRHX2AD
MACRO SDFFNSRHX4AD
    CLASS CORE ;
    FOREIGN SDFFNSRHX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 1.110 5.265 1.375 ;
        END
        AntennaGateArea 0.194 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.985 0.860 3.335 1.050 ;
        END
        AntennaGateArea 0.077 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 0.860 3.810 1.340 ;
        RECT  2.860 1.190 3.550 1.340 ;
        END
        AntennaGateArea 0.125 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.720 0.960 11.840 1.220 ;
        RECT  10.195 1.100 11.720 1.220 ;
        RECT  9.685 1.100 10.195 1.330 ;
        RECT  9.085 1.100 9.685 1.220 ;
        RECT  8.965 0.910 9.085 1.220 ;
        END
        AntennaGateArea 0.226 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.115 1.730 13.255 1.850 ;
        RECT  12.995 0.910 13.115 1.850 ;
        RECT  12.950 0.910 12.995 1.515 ;
        RECT  12.670 0.910 12.950 1.030 ;
        END
        AntennaDiffArea 0.198 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.395 1.005 14.490 1.515 ;
        RECT  14.225 0.365 14.395 2.175 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.920 2.260 1.375 ;
        END
        AntennaGateArea 0.144 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.110 0.770 1.375 ;
        END
        AntennaGateArea 0.167 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.755 -0.210 14.840 0.210 ;
        RECT  14.585 -0.210 14.755 0.795 ;
        RECT  14.010 -0.210 14.585 0.210 ;
        RECT  13.750 -0.210 14.010 0.310 ;
        RECT  13.330 -0.210 13.750 0.210 ;
        RECT  13.070 -0.210 13.330 0.310 ;
        RECT  12.460 -0.210 13.070 0.210 ;
        RECT  12.200 -0.210 12.460 0.310 ;
        RECT  10.210 -0.210 12.200 0.210 ;
        RECT  10.040 -0.210 10.210 0.260 ;
        RECT  8.940 -0.210 10.040 0.210 ;
        RECT  8.770 -0.210 8.940 0.260 ;
        RECT  8.130 -0.210 8.770 0.210 ;
        RECT  7.870 -0.210 8.130 0.230 ;
        RECT  7.240 -0.210 7.870 0.210 ;
        RECT  6.980 -0.210 7.240 0.230 ;
        RECT  5.280 -0.210 6.980 0.210 ;
        RECT  4.760 -0.210 5.280 0.230 ;
        RECT  4.210 -0.210 4.760 0.210 ;
        RECT  3.690 -0.210 4.210 0.230 ;
        RECT  1.895 -0.210 3.690 0.210 ;
        RECT  1.725 -0.210 1.895 0.450 ;
        RECT  0.610 -0.210 1.725 0.210 ;
        RECT  0.470 -0.210 0.610 0.750 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.755 2.310 14.840 2.730 ;
        RECT  14.585 1.635 14.755 2.730 ;
        RECT  14.035 2.310 14.585 2.730 ;
        RECT  13.865 1.960 14.035 2.730 ;
        RECT  13.655 2.310 13.865 2.730 ;
        RECT  13.395 2.210 13.655 2.730 ;
        RECT  11.980 2.310 13.395 2.730 ;
        RECT  11.720 2.220 11.980 2.730 ;
        RECT  9.340 2.310 11.720 2.730 ;
        RECT  9.170 2.260 9.340 2.730 ;
        RECT  8.410 2.310 9.170 2.730 ;
        RECT  8.240 2.260 8.410 2.730 ;
        RECT  6.945 2.310 8.240 2.730 ;
        RECT  6.775 2.260 6.945 2.730 ;
        RECT  5.300 2.310 6.775 2.730 ;
        RECT  4.780 2.260 5.300 2.730 ;
        RECT  4.280 2.310 4.780 2.730 ;
        RECT  3.760 2.260 4.280 2.730 ;
        RECT  2.605 2.310 3.760 2.730 ;
        RECT  2.345 2.290 2.605 2.730 ;
        RECT  1.510 2.310 2.345 2.730 ;
        RECT  1.250 2.265 1.510 2.730 ;
        RECT  0.575 2.310 1.250 2.730 ;
        RECT  0.405 2.105 0.575 2.730 ;
        RECT  0.000 2.310 0.405 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 14.840 2.520 ;
        LAYER M1 ;
        RECT  13.905 1.015 14.080 1.275 ;
        RECT  13.785 0.430 13.905 1.840 ;
        RECT  12.800 0.430 13.785 0.550 ;
        RECT  13.700 1.015 13.785 1.275 ;
        RECT  13.500 1.720 13.785 1.840 ;
        RECT  13.545 1.420 13.655 1.590 ;
        RECT  13.545 0.670 13.635 0.905 ;
        RECT  13.425 0.670 13.545 1.590 ;
        RECT  13.380 1.720 13.500 2.090 ;
        RECT  12.325 0.670 13.425 0.790 ;
        RECT  13.235 1.125 13.425 1.295 ;
        RECT  12.855 1.970 13.380 2.090 ;
        RECT  12.685 1.795 12.855 2.090 ;
        RECT  12.690 1.490 12.830 1.610 ;
        RECT  12.630 0.355 12.800 0.550 ;
        RECT  12.570 1.190 12.690 1.610 ;
        RECT  11.570 1.970 12.685 2.090 ;
        RECT  11.755 0.430 12.630 0.550 ;
        RECT  12.085 1.190 12.570 1.310 ;
        RECT  11.330 1.430 12.450 1.550 ;
        RECT  12.205 0.670 12.325 0.975 ;
        RECT  11.965 0.670 12.085 1.310 ;
        RECT  11.535 0.670 11.965 0.790 ;
        RECT  11.635 0.380 11.755 0.550 ;
        RECT  10.450 0.380 11.635 0.500 ;
        RECT  11.480 1.970 11.570 2.115 ;
        RECT  11.415 0.620 11.535 0.790 ;
        RECT  10.355 1.995 11.480 2.115 ;
        RECT  10.060 0.620 11.415 0.740 ;
        RECT  11.205 1.430 11.330 1.875 ;
        RECT  7.980 1.755 11.205 1.875 ;
        RECT  9.625 0.860 11.100 0.980 ;
        RECT  8.655 1.515 10.995 1.635 ;
        RECT  9.940 0.380 10.060 0.740 ;
        RECT  9.785 2.020 10.045 2.190 ;
        RECT  2.135 0.380 9.940 0.500 ;
        RECT  7.855 2.020 9.785 2.140 ;
        RECT  9.505 0.620 9.625 0.980 ;
        RECT  9.365 0.620 9.505 0.790 ;
        RECT  8.655 0.670 9.365 0.790 ;
        RECT  8.535 0.670 8.655 1.635 ;
        RECT  8.100 1.410 8.535 1.530 ;
        RECT  8.295 0.635 8.415 1.285 ;
        RECT  4.920 0.635 8.295 0.755 ;
        RECT  7.980 1.165 8.295 1.285 ;
        RECT  7.740 0.925 8.125 1.045 ;
        RECT  7.860 1.165 7.980 1.875 ;
        RECT  7.595 2.020 7.855 2.190 ;
        RECT  7.620 0.925 7.740 1.870 ;
        RECT  7.060 0.925 7.620 1.045 ;
        RECT  6.075 1.750 7.620 1.870 ;
        RECT  5.825 2.020 7.595 2.140 ;
        RECT  7.325 1.340 7.445 1.600 ;
        RECT  6.455 1.480 7.325 1.600 ;
        RECT  6.930 0.905 7.060 1.045 ;
        RECT  6.290 0.905 6.930 1.025 ;
        RECT  5.825 1.160 6.790 1.280 ;
        RECT  6.195 1.410 6.455 1.600 ;
        RECT  6.030 0.880 6.290 1.025 ;
        RECT  5.710 1.160 5.825 2.140 ;
        RECT  5.705 1.070 5.710 2.140 ;
        RECT  5.590 1.070 5.705 1.330 ;
        RECT  1.820 2.020 5.705 2.140 ;
        RECT  4.535 1.780 5.560 1.900 ;
        RECT  4.800 0.635 4.920 1.620 ;
        RECT  4.655 1.500 4.800 1.620 ;
        RECT  4.550 0.620 4.670 1.230 ;
        RECT  4.050 0.620 4.550 0.740 ;
        RECT  4.535 1.105 4.550 1.230 ;
        RECT  4.415 1.105 4.535 1.900 ;
        RECT  4.295 0.860 4.430 0.980 ;
        RECT  4.170 0.860 4.295 1.900 ;
        RECT  2.780 1.780 4.170 1.900 ;
        RECT  3.930 0.620 4.050 1.650 ;
        RECT  2.795 0.620 3.930 0.740 ;
        RECT  2.900 1.530 3.930 1.650 ;
        RECT  2.740 1.515 2.780 1.900 ;
        RECT  2.660 0.855 2.740 1.900 ;
        RECT  2.620 0.855 2.660 1.635 ;
        RECT  2.500 1.730 2.540 1.900 ;
        RECT  2.500 0.670 2.515 0.790 ;
        RECT  2.380 0.670 2.500 1.900 ;
        RECT  2.255 0.670 2.380 0.790 ;
        RECT  2.340 1.730 2.380 1.900 ;
        RECT  2.015 0.380 2.135 0.690 ;
        RECT  1.090 0.570 2.015 0.690 ;
        RECT  1.700 1.135 1.820 2.140 ;
        RECT  1.520 1.135 1.700 1.255 ;
        RECT  1.400 0.815 1.520 1.255 ;
        RECT  1.260 0.815 1.400 0.935 ;
        RECT  1.350 1.135 1.400 1.255 ;
        RECT  1.230 1.135 1.350 1.395 ;
        RECT  0.850 0.330 1.250 0.450 ;
        RECT  1.090 1.575 1.205 2.005 ;
        RECT  0.970 0.570 1.090 2.005 ;
        RECT  0.730 0.330 0.850 0.990 ;
        RECT  0.265 0.870 0.730 0.990 ;
        RECT  0.215 0.635 0.265 0.990 ;
        RECT  0.215 1.565 0.265 1.735 ;
        RECT  0.095 0.635 0.215 1.735 ;
    END
END SDFFNSRHX4AD
MACRO SDFFNSRHX8AD
    CLASS CORE ;
    FOREIGN SDFFNSRHX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 1.110 5.265 1.375 ;
        END
        AntennaGateArea 0.235 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.985 0.860 3.335 1.050 ;
        END
        AntennaGateArea 0.101 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 0.860 3.810 1.340 ;
        RECT  2.860 1.190 3.550 1.340 ;
        END
        AntennaGateArea 0.149 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.720 0.960 11.840 1.220 ;
        RECT  10.195 1.100 11.720 1.220 ;
        RECT  9.685 1.100 10.195 1.330 ;
        RECT  9.085 1.100 9.685 1.220 ;
        RECT  8.965 0.910 9.085 1.220 ;
        END
        AntennaGateArea 0.237 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.995 0.910 13.255 1.850 ;
        RECT  12.810 0.910 12.995 1.515 ;
        RECT  12.670 0.910 12.810 1.030 ;
        END
        AntennaDiffArea 0.204 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.065 0.365 15.235 2.175 ;
        RECT  14.515 1.005 15.065 1.515 ;
        RECT  14.345 0.365 14.515 2.175 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.930 2.260 1.375 ;
        END
        AntennaGateArea 0.144 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.110 0.770 1.375 ;
        END
        AntennaGateArea 0.255 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.595 -0.210 15.680 0.210 ;
        RECT  15.425 -0.210 15.595 0.795 ;
        RECT  14.875 -0.210 15.425 0.210 ;
        RECT  14.705 -0.210 14.875 0.795 ;
        RECT  14.130 -0.210 14.705 0.210 ;
        RECT  13.870 -0.210 14.130 0.310 ;
        RECT  13.330 -0.210 13.870 0.210 ;
        RECT  13.070 -0.210 13.330 0.310 ;
        RECT  12.460 -0.210 13.070 0.210 ;
        RECT  12.200 -0.210 12.460 0.310 ;
        RECT  10.260 -0.210 12.200 0.210 ;
        RECT  10.090 -0.210 10.260 0.260 ;
        RECT  8.890 -0.210 10.090 0.210 ;
        RECT  8.720 -0.210 8.890 0.260 ;
        RECT  8.085 -0.210 8.720 0.210 ;
        RECT  7.915 -0.210 8.085 0.260 ;
        RECT  7.195 -0.210 7.915 0.210 ;
        RECT  7.025 -0.210 7.195 0.255 ;
        RECT  5.280 -0.210 7.025 0.210 ;
        RECT  4.760 -0.210 5.280 0.260 ;
        RECT  4.210 -0.210 4.760 0.210 ;
        RECT  3.690 -0.210 4.210 0.260 ;
        RECT  1.895 -0.210 3.690 0.210 ;
        RECT  1.725 -0.210 1.895 0.450 ;
        RECT  0.610 -0.210 1.725 0.210 ;
        RECT  0.470 -0.210 0.610 0.750 ;
        RECT  0.000 -0.210 0.470 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.595 2.310 15.680 2.730 ;
        RECT  15.425 1.485 15.595 2.730 ;
        RECT  14.875 2.310 15.425 2.730 ;
        RECT  14.705 1.635 14.875 2.730 ;
        RECT  14.155 2.310 14.705 2.730 ;
        RECT  13.985 1.960 14.155 2.730 ;
        RECT  13.655 2.310 13.985 2.730 ;
        RECT  13.395 2.210 13.655 2.730 ;
        RECT  11.980 2.310 13.395 2.730 ;
        RECT  11.720 2.220 11.980 2.730 ;
        RECT  9.390 2.310 11.720 2.730 ;
        RECT  9.220 2.260 9.390 2.730 ;
        RECT  8.410 2.310 9.220 2.730 ;
        RECT  8.240 2.260 8.410 2.730 ;
        RECT  6.945 2.310 8.240 2.730 ;
        RECT  6.775 2.260 6.945 2.730 ;
        RECT  5.300 2.310 6.775 2.730 ;
        RECT  4.780 2.260 5.300 2.730 ;
        RECT  4.280 2.310 4.780 2.730 ;
        RECT  3.760 2.260 4.280 2.730 ;
        RECT  2.560 2.310 3.760 2.730 ;
        RECT  2.390 2.265 2.560 2.730 ;
        RECT  1.465 2.310 2.390 2.730 ;
        RECT  1.295 2.175 1.465 2.730 ;
        RECT  0.565 2.310 1.295 2.730 ;
        RECT  0.395 2.265 0.565 2.730 ;
        RECT  0.000 2.310 0.395 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 15.680 2.520 ;
        LAYER M1 ;
        RECT  14.025 1.015 14.200 1.275 ;
        RECT  13.905 0.430 14.025 1.840 ;
        RECT  12.800 0.430 13.905 0.550 ;
        RECT  13.820 1.015 13.905 1.275 ;
        RECT  13.500 1.720 13.905 1.840 ;
        RECT  13.640 0.735 13.755 0.905 ;
        RECT  13.640 1.420 13.755 1.590 ;
        RECT  13.520 0.670 13.640 1.590 ;
        RECT  12.325 0.670 13.520 0.790 ;
        RECT  13.375 1.055 13.520 1.225 ;
        RECT  13.380 1.720 13.500 2.090 ;
        RECT  12.855 1.970 13.380 2.090 ;
        RECT  12.685 1.890 12.855 2.090 ;
        RECT  12.690 1.635 12.830 1.755 ;
        RECT  12.630 0.330 12.800 0.550 ;
        RECT  12.570 1.190 12.690 1.755 ;
        RECT  11.570 1.970 12.685 2.090 ;
        RECT  11.755 0.430 12.630 0.550 ;
        RECT  12.085 1.190 12.570 1.310 ;
        RECT  11.240 1.430 12.450 1.550 ;
        RECT  12.205 0.670 12.325 0.975 ;
        RECT  11.965 0.670 12.085 1.310 ;
        RECT  11.535 0.670 11.965 0.790 ;
        RECT  11.635 0.380 11.755 0.550 ;
        RECT  10.450 0.380 11.635 0.500 ;
        RECT  11.480 1.970 11.570 2.115 ;
        RECT  11.415 0.620 11.535 0.790 ;
        RECT  10.355 1.995 11.480 2.115 ;
        RECT  10.060 0.620 11.415 0.740 ;
        RECT  11.115 1.430 11.240 1.875 ;
        RECT  9.685 1.755 11.115 1.875 ;
        RECT  9.625 0.860 11.100 0.980 ;
        RECT  8.655 1.515 10.995 1.635 ;
        RECT  9.940 0.380 10.060 0.740 ;
        RECT  9.785 2.020 10.045 2.190 ;
        RECT  7.545 0.380 9.940 0.500 ;
        RECT  7.845 2.020 9.785 2.140 ;
        RECT  9.425 1.755 9.685 1.900 ;
        RECT  9.505 0.620 9.625 0.980 ;
        RECT  9.365 0.620 9.505 0.790 ;
        RECT  7.980 1.755 9.425 1.875 ;
        RECT  8.655 0.670 9.365 0.790 ;
        RECT  8.535 0.670 8.655 1.635 ;
        RECT  8.100 1.410 8.535 1.530 ;
        RECT  8.295 0.635 8.415 1.285 ;
        RECT  4.920 0.635 8.295 0.755 ;
        RECT  7.980 1.165 8.295 1.285 ;
        RECT  7.740 0.925 8.125 1.045 ;
        RECT  7.860 1.165 7.980 1.875 ;
        RECT  7.585 2.020 7.845 2.190 ;
        RECT  7.620 0.925 7.740 1.870 ;
        RECT  7.060 0.925 7.620 1.045 ;
        RECT  6.075 1.750 7.620 1.870 ;
        RECT  5.825 2.020 7.585 2.140 ;
        RECT  7.285 0.345 7.545 0.500 ;
        RECT  7.325 1.340 7.445 1.600 ;
        RECT  6.455 1.480 7.325 1.600 ;
        RECT  2.135 0.380 7.285 0.500 ;
        RECT  6.930 0.905 7.060 1.045 ;
        RECT  6.290 0.905 6.930 1.025 ;
        RECT  5.825 1.160 6.790 1.280 ;
        RECT  6.195 1.410 6.455 1.600 ;
        RECT  6.030 0.880 6.290 1.025 ;
        RECT  5.710 1.160 5.825 2.140 ;
        RECT  5.705 1.070 5.710 2.140 ;
        RECT  5.590 1.070 5.705 1.330 ;
        RECT  1.820 2.020 5.705 2.140 ;
        RECT  4.535 1.780 5.560 1.900 ;
        RECT  4.800 0.635 4.920 1.620 ;
        RECT  4.655 1.500 4.800 1.620 ;
        RECT  4.550 0.620 4.670 1.230 ;
        RECT  4.050 0.620 4.550 0.740 ;
        RECT  4.535 1.105 4.550 1.230 ;
        RECT  4.415 1.105 4.535 1.900 ;
        RECT  4.295 0.860 4.430 0.980 ;
        RECT  4.170 0.860 4.295 1.900 ;
        RECT  2.780 1.780 4.170 1.900 ;
        RECT  3.930 0.620 4.050 1.650 ;
        RECT  2.780 0.620 3.930 0.740 ;
        RECT  2.900 1.530 3.930 1.650 ;
        RECT  2.740 1.515 2.780 1.900 ;
        RECT  2.660 0.855 2.740 1.900 ;
        RECT  2.620 0.855 2.660 1.635 ;
        RECT  2.500 1.730 2.540 1.900 ;
        RECT  2.380 0.645 2.500 1.900 ;
        RECT  2.300 0.645 2.380 0.815 ;
        RECT  2.340 1.730 2.380 1.900 ;
        RECT  2.015 0.380 2.135 0.690 ;
        RECT  1.090 0.570 2.015 0.690 ;
        RECT  1.700 1.115 1.820 2.140 ;
        RECT  1.520 1.115 1.700 1.255 ;
        RECT  1.400 0.815 1.520 1.255 ;
        RECT  1.260 0.815 1.400 0.935 ;
        RECT  1.350 1.115 1.400 1.255 ;
        RECT  1.230 1.115 1.350 1.375 ;
        RECT  0.850 0.330 1.250 0.450 ;
        RECT  1.090 1.575 1.205 2.005 ;
        RECT  0.970 0.570 1.090 2.005 ;
        RECT  0.730 0.330 0.850 0.990 ;
        RECT  0.250 0.870 0.730 0.990 ;
        RECT  0.215 0.330 0.250 0.990 ;
        RECT  0.215 1.435 0.245 1.955 ;
        RECT  0.095 0.330 0.215 1.955 ;
    END
END SDFFNSRHX8AD
MACRO SDFFQX1AD
    CLASS CORE ;
    FOREIGN SDFFQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.015 1.080 1.275 ;
        RECT  0.910 1.015 1.050 1.375 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.430 1.470 1.550 ;
        RECT  1.200 1.430 1.320 1.770 ;
        RECT  0.210 1.650 1.200 1.770 ;
        RECT  0.210 1.005 0.485 1.265 ;
        RECT  0.070 1.005 0.210 1.770 ;
        END
        AntennaGateArea 0.119 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.790 0.380 6.930 2.085 ;
        RECT  6.735 0.380 6.790 0.550 ;
        RECT  6.760 1.565 6.790 2.085 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.390 0.910 1.740 1.115 ;
        END
        AntennaGateArea 0.071 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.225 1.380 3.615 1.620 ;
        RECT  3.105 1.020 3.225 1.620 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.545 -0.210 7.000 0.210 ;
        RECT  6.375 -0.210 6.545 0.500 ;
        RECT  6.025 -0.210 6.375 0.210 ;
        RECT  5.765 -0.210 6.025 0.770 ;
        RECT  4.755 -0.210 5.765 0.210 ;
        RECT  4.495 -0.210 4.755 0.430 ;
        RECT  3.615 -0.210 4.495 0.210 ;
        RECT  3.355 -0.210 3.615 0.420 ;
        RECT  2.950 -0.210 3.355 0.210 ;
        RECT  2.690 -0.210 2.950 0.420 ;
        RECT  1.300 -0.210 2.690 0.210 ;
        RECT  1.040 -0.210 1.300 0.300 ;
        RECT  0.265 -0.210 1.040 0.210 ;
        RECT  0.095 -0.210 0.265 0.495 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.590 2.310 7.000 2.730 ;
        RECT  6.330 2.010 6.590 2.730 ;
        RECT  5.930 2.310 6.330 2.730 ;
        RECT  5.670 2.025 5.930 2.730 ;
        RECT  4.755 2.310 5.670 2.730 ;
        RECT  4.495 2.220 4.755 2.730 ;
        RECT  3.715 2.310 4.495 2.730 ;
        RECT  3.455 2.220 3.715 2.730 ;
        RECT  2.995 2.310 3.455 2.730 ;
        RECT  2.735 2.220 2.995 2.730 ;
        RECT  1.320 2.310 2.735 2.730 ;
        RECT  1.060 2.220 1.320 2.730 ;
        RECT  0.255 2.310 1.060 2.730 ;
        RECT  0.085 1.890 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.550 0.780 6.670 1.445 ;
        RECT  6.395 0.780 6.550 0.900 ;
        RECT  6.265 1.325 6.550 1.445 ;
        RECT  6.120 1.085 6.430 1.205 ;
        RECT  6.225 0.730 6.395 0.900 ;
        RECT  6.095 1.325 6.265 1.750 ;
        RECT  6.000 0.975 6.120 1.205 ;
        RECT  5.850 1.325 6.095 1.445 ;
        RECT  5.365 0.975 6.000 1.095 ;
        RECT  5.590 1.275 5.850 1.445 ;
        RECT  5.270 0.330 5.530 0.500 ;
        RECT  5.195 0.625 5.365 1.780 ;
        RECT  5.075 0.380 5.270 0.500 ;
        RECT  5.075 2.070 5.265 2.190 ;
        RECT  4.955 0.380 5.075 2.190 ;
        RECT  4.555 0.620 4.955 0.740 ;
        RECT  4.930 1.980 4.955 2.190 ;
        RECT  2.600 1.980 4.930 2.100 ;
        RECT  4.705 1.045 4.825 1.860 ;
        RECT  3.975 1.740 4.705 1.860 ;
        RECT  4.435 0.620 4.555 1.310 ;
        RECT  4.335 1.050 4.435 1.310 ;
        RECT  4.215 1.495 4.375 1.615 ;
        RECT  4.215 0.455 4.305 0.920 ;
        RECT  4.095 0.330 4.215 1.615 ;
        RECT  3.835 0.330 4.095 0.590 ;
        RECT  3.855 0.755 3.975 1.860 ;
        RECT  3.685 0.755 3.855 0.875 ;
        RECT  2.840 1.740 3.855 1.860 ;
        RECT  3.595 1.000 3.715 1.260 ;
        RECT  3.505 1.000 3.595 1.120 ;
        RECT  3.385 0.540 3.505 1.120 ;
        RECT  2.360 0.540 3.385 0.660 ;
        RECT  2.600 0.780 3.255 0.900 ;
        RECT  2.720 1.260 2.840 1.860 ;
        RECT  2.480 0.780 2.600 2.190 ;
        RECT  2.290 2.020 2.480 2.190 ;
        RECT  2.240 0.540 2.360 1.900 ;
        RECT  2.120 2.020 2.290 2.140 ;
        RECT  2.060 0.540 2.240 0.730 ;
        RECT  2.000 0.920 2.120 2.140 ;
        RECT  1.860 0.920 2.000 1.040 ;
        RECT  1.670 0.380 1.930 0.540 ;
        RECT  1.760 1.640 1.880 2.160 ;
        RECT  0.690 1.980 1.760 2.100 ;
        RECT  0.670 0.420 1.670 0.540 ;
        RECT  0.745 0.660 1.440 0.780 ;
        RECT  0.745 1.270 0.780 1.530 ;
        RECT  0.625 0.660 0.745 1.530 ;
        RECT  0.430 1.890 0.690 2.100 ;
        RECT  0.410 0.380 0.670 0.540 ;
        RECT  0.330 0.660 0.625 0.880 ;
        RECT  0.330 1.410 0.625 1.530 ;
    END
END SDFFQX1AD
MACRO SDFFQX2AD
    CLASS CORE ;
    FOREIGN SDFFQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.190 1.655 1.330 ;
        RECT  0.900 1.170 1.160 1.330 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.450 1.470 1.610 ;
        RECT  1.200 1.450 1.320 1.770 ;
        RECT  0.210 1.650 1.200 1.770 ;
        RECT  0.210 1.005 0.485 1.265 ;
        RECT  0.070 1.005 0.210 1.770 ;
        END
        AntennaGateArea 0.119 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.770 0.360 6.930 2.180 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.480 0.910 1.740 1.070 ;
        RECT  0.865 0.910 1.480 1.050 ;
        END
        AntennaGateArea 0.071 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.225 1.380 3.615 1.620 ;
        RECT  3.105 1.020 3.225 1.620 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.560 -0.210 7.000 0.210 ;
        RECT  6.340 -0.210 6.560 0.445 ;
        RECT  6.025 -0.210 6.340 0.210 ;
        RECT  5.765 -0.210 6.025 0.330 ;
        RECT  4.675 -0.210 5.765 0.210 ;
        RECT  4.415 -0.210 4.675 0.630 ;
        RECT  3.615 -0.210 4.415 0.210 ;
        RECT  3.355 -0.210 3.615 0.420 ;
        RECT  2.950 -0.210 3.355 0.210 ;
        RECT  2.690 -0.210 2.950 0.420 ;
        RECT  1.300 -0.210 2.690 0.210 ;
        RECT  1.040 -0.210 1.300 0.300 ;
        RECT  0.265 -0.210 1.040 0.210 ;
        RECT  0.095 -0.210 0.265 0.495 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.555 2.310 7.000 2.730 ;
        RECT  6.385 2.060 6.555 2.730 ;
        RECT  5.905 2.310 6.385 2.730 ;
        RECT  5.685 2.075 5.905 2.730 ;
        RECT  4.645 2.310 5.685 2.730 ;
        RECT  4.385 2.220 4.645 2.730 ;
        RECT  3.715 2.310 4.385 2.730 ;
        RECT  3.455 2.220 3.715 2.730 ;
        RECT  2.995 2.310 3.455 2.730 ;
        RECT  2.735 2.220 2.995 2.730 ;
        RECT  1.320 2.310 2.735 2.730 ;
        RECT  1.060 2.220 1.320 2.730 ;
        RECT  0.255 2.310 1.060 2.730 ;
        RECT  0.085 1.890 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.530 0.780 6.650 1.490 ;
        RECT  6.270 0.780 6.530 0.900 ;
        RECT  6.270 1.370 6.530 1.490 ;
        RECT  6.040 1.060 6.410 1.230 ;
        RECT  6.145 0.625 6.270 0.900 ;
        RECT  6.100 1.370 6.270 1.750 ;
        RECT  6.100 0.625 6.145 0.795 ;
        RECT  5.765 1.370 6.100 1.490 ;
        RECT  5.920 0.975 6.040 1.230 ;
        RECT  5.285 0.975 5.920 1.095 ;
        RECT  5.505 1.275 5.765 1.490 ;
        RECT  5.255 0.330 5.515 0.500 ;
        RECT  5.235 0.625 5.285 1.095 ;
        RECT  4.995 0.380 5.255 0.500 ;
        RECT  5.115 0.625 5.235 1.780 ;
        RECT  4.995 2.070 5.155 2.190 ;
        RECT  4.875 0.380 4.995 2.190 ;
        RECT  4.455 0.750 4.875 0.870 ;
        RECT  2.600 1.980 4.875 2.100 ;
        RECT  4.635 1.020 4.755 1.860 ;
        RECT  3.975 1.740 4.635 1.860 ;
        RECT  4.335 0.750 4.455 1.290 ;
        RECT  4.215 1.465 4.355 1.585 ;
        RECT  4.095 0.375 4.215 1.585 ;
        RECT  3.900 0.375 4.095 0.545 ;
        RECT  3.855 0.755 3.975 1.860 ;
        RECT  3.685 0.755 3.855 0.875 ;
        RECT  2.840 1.740 3.855 1.860 ;
        RECT  3.595 1.000 3.715 1.260 ;
        RECT  3.505 1.000 3.595 1.120 ;
        RECT  3.385 0.540 3.505 1.120 ;
        RECT  2.360 0.540 3.385 0.660 ;
        RECT  2.600 0.780 3.255 0.900 ;
        RECT  2.720 1.260 2.840 1.860 ;
        RECT  2.480 0.780 2.600 2.190 ;
        RECT  2.290 2.020 2.480 2.190 ;
        RECT  2.240 0.540 2.360 1.900 ;
        RECT  2.120 2.020 2.290 2.140 ;
        RECT  2.060 0.540 2.240 0.730 ;
        RECT  2.000 0.920 2.120 2.140 ;
        RECT  1.860 0.920 2.000 1.040 ;
        RECT  1.670 0.380 1.930 0.540 ;
        RECT  1.760 1.640 1.880 2.160 ;
        RECT  0.690 1.980 1.760 2.100 ;
        RECT  0.670 0.420 1.670 0.540 ;
        RECT  0.745 0.660 1.440 0.780 ;
        RECT  0.745 1.270 0.780 1.530 ;
        RECT  0.625 0.660 0.745 1.530 ;
        RECT  0.430 1.890 0.690 2.100 ;
        RECT  0.410 0.380 0.670 0.540 ;
        RECT  0.330 0.660 0.625 0.880 ;
        RECT  0.330 1.410 0.625 1.530 ;
    END
END SDFFQX2AD
MACRO SDFFQX4AD
    CLASS CORE ;
    FOREIGN SDFFQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 1.190 1.375 1.330 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.470 1.665 1.610 ;
        RECT  1.210 1.470 1.470 1.760 ;
        RECT  0.200 1.640 1.210 1.760 ;
        RECT  0.200 1.005 0.320 1.265 ;
        RECT  0.080 1.005 0.200 1.760 ;
        END
        AntennaGateArea 0.119 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.065 0.365 8.235 2.115 ;
        RECT  7.910 1.005 8.065 1.515 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.980 1.890 1.375 ;
        RECT  1.635 0.980 1.750 1.350 ;
        RECT  1.530 1.230 1.635 1.350 ;
        END
        AntennaGateArea 0.071 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.825 1.430 3.335 1.610 ;
        END
        AntennaGateArea 0.091 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.595 -0.210 8.680 0.210 ;
        RECT  8.425 -0.210 8.595 0.795 ;
        RECT  7.875 -0.210 8.425 0.210 ;
        RECT  7.705 -0.210 7.875 0.535 ;
        RECT  7.240 -0.210 7.705 0.210 ;
        RECT  6.980 -0.210 7.240 0.435 ;
        RECT  5.700 -0.210 6.980 0.210 ;
        RECT  5.440 -0.210 5.700 0.505 ;
        RECT  4.165 -0.210 5.440 0.210 ;
        RECT  3.995 -0.210 4.165 0.550 ;
        RECT  3.090 -0.210 3.995 0.210 ;
        RECT  2.830 -0.210 3.090 0.540 ;
        RECT  1.330 -0.210 2.830 0.210 ;
        RECT  1.070 -0.210 1.330 0.290 ;
        RECT  0.230 -0.210 1.070 0.210 ;
        RECT  0.110 -0.210 0.230 0.520 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.595 2.310 8.680 2.730 ;
        RECT  8.425 1.425 8.595 2.730 ;
        RECT  7.875 2.310 8.425 2.730 ;
        RECT  7.705 1.765 7.875 2.730 ;
        RECT  7.145 2.310 7.705 2.730 ;
        RECT  6.975 1.945 7.145 2.730 ;
        RECT  5.760 2.310 6.975 2.730 ;
        RECT  5.640 1.505 5.760 2.730 ;
        RECT  4.810 2.310 5.640 2.730 ;
        RECT  4.550 2.220 4.810 2.730 ;
        RECT  3.790 2.310 4.550 2.730 ;
        RECT  3.530 2.220 3.790 2.730 ;
        RECT  3.070 2.310 3.530 2.730 ;
        RECT  2.810 2.220 3.070 2.730 ;
        RECT  1.330 2.310 2.810 2.730 ;
        RECT  1.070 2.120 1.330 2.730 ;
        RECT  0.255 2.310 1.070 2.730 ;
        RECT  0.085 1.890 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.680 2.520 ;
        LAYER M1 ;
        RECT  7.670 0.720 7.790 1.615 ;
        RECT  7.365 0.720 7.670 0.890 ;
        RECT  6.830 1.495 7.670 1.615 ;
        RECT  7.200 1.020 7.550 1.280 ;
        RECT  7.080 0.625 7.200 1.375 ;
        RECT  4.810 0.625 7.080 0.745 ;
        RECT  6.450 1.255 7.080 1.375 ;
        RECT  6.710 1.495 6.830 2.120 ;
        RECT  5.210 0.910 6.730 1.030 ;
        RECT  6.250 1.255 6.450 2.075 ;
        RECT  5.520 1.255 6.250 1.375 ;
        RECT  5.400 1.255 5.520 2.050 ;
        RECT  5.090 1.930 5.400 2.050 ;
        RECT  5.090 0.910 5.210 1.810 ;
        RECT  4.520 0.910 5.090 1.030 ;
        RECT  4.850 1.690 5.090 1.810 ;
        RECT  4.970 1.930 5.090 2.190 ;
        RECT  4.855 1.150 4.970 1.270 ;
        RECT  4.710 1.150 4.855 1.570 ;
        RECT  4.730 1.690 4.850 2.100 ;
        RECT  3.340 1.980 4.730 2.100 ;
        RECT  4.610 1.450 4.710 1.570 ;
        RECT  4.495 0.330 4.665 0.790 ;
        RECT  4.490 1.450 4.610 1.860 ;
        RECT  4.400 0.910 4.520 1.220 ;
        RECT  4.280 0.670 4.495 0.790 ;
        RECT  4.010 1.740 4.490 1.860 ;
        RECT  4.280 1.355 4.370 1.615 ;
        RECT  4.160 0.670 4.280 1.615 ;
        RECT  3.890 0.675 4.010 1.860 ;
        RECT  3.785 0.675 3.890 0.805 ;
        RECT  3.810 1.190 3.890 1.860 ;
        RECT  2.640 1.190 3.810 1.310 ;
        RECT  3.615 0.635 3.785 0.805 ;
        RECT  2.390 0.950 3.770 1.070 ;
        RECT  2.630 0.710 3.470 0.830 ;
        RECT  3.220 1.730 3.340 2.100 ;
        RECT  2.665 1.980 3.220 2.100 ;
        RECT  2.590 1.980 2.665 2.140 ;
        RECT  2.510 0.380 2.630 0.830 ;
        RECT  2.545 1.980 2.590 2.190 ;
        RECT  2.330 2.020 2.545 2.190 ;
        RECT  2.130 0.380 2.510 0.500 ;
        RECT  2.250 0.640 2.390 1.875 ;
        RECT  2.130 2.020 2.330 2.140 ;
        RECT  2.010 0.380 2.130 2.140 ;
        RECT  1.770 0.495 1.890 0.790 ;
        RECT  1.770 1.880 1.890 2.145 ;
        RECT  0.655 0.495 1.770 0.615 ;
        RECT  0.440 1.880 1.770 2.000 ;
        RECT  1.170 0.760 1.430 1.005 ;
        RECT  0.560 0.760 1.170 0.880 ;
        RECT  0.560 1.400 0.850 1.520 ;
        RECT  0.485 0.395 0.655 0.615 ;
        RECT  0.440 0.760 0.560 1.520 ;
        RECT  0.330 0.760 0.440 0.880 ;
        RECT  0.330 1.400 0.440 1.520 ;
    END
END SDFFQX4AD
MACRO SDFFQXLAD
    CLASS CORE ;
    FOREIGN SDFFQXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.015 1.080 1.275 ;
        RECT  0.910 1.015 1.050 1.375 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.430 1.470 1.550 ;
        RECT  1.200 1.430 1.320 1.770 ;
        RECT  0.210 1.650 1.200 1.770 ;
        RECT  0.210 1.005 0.485 1.265 ;
        RECT  0.070 1.005 0.210 1.770 ;
        END
        AntennaGateArea 0.119 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.790 0.390 6.930 2.085 ;
        RECT  6.735 0.390 6.790 0.560 ;
        RECT  6.760 1.825 6.790 2.085 ;
        END
        AntennaDiffArea 0.138 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.390 0.910 1.740 1.115 ;
        END
        AntennaGateArea 0.071 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.225 1.380 3.615 1.620 ;
        RECT  3.105 1.020 3.225 1.620 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.545 -0.210 7.000 0.210 ;
        RECT  6.375 -0.210 6.545 0.560 ;
        RECT  6.025 -0.210 6.375 0.210 ;
        RECT  5.765 -0.210 6.025 0.770 ;
        RECT  4.755 -0.210 5.765 0.210 ;
        RECT  4.495 -0.210 4.755 0.430 ;
        RECT  3.615 -0.210 4.495 0.210 ;
        RECT  3.355 -0.210 3.615 0.420 ;
        RECT  2.950 -0.210 3.355 0.210 ;
        RECT  2.690 -0.210 2.950 0.420 ;
        RECT  1.300 -0.210 2.690 0.210 ;
        RECT  1.040 -0.210 1.300 0.300 ;
        RECT  0.265 -0.210 1.040 0.210 ;
        RECT  0.095 -0.210 0.265 0.495 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.590 2.310 7.000 2.730 ;
        RECT  6.330 2.010 6.590 2.730 ;
        RECT  5.930 2.310 6.330 2.730 ;
        RECT  5.670 2.025 5.930 2.730 ;
        RECT  4.755 2.310 5.670 2.730 ;
        RECT  4.495 2.220 4.755 2.730 ;
        RECT  3.715 2.310 4.495 2.730 ;
        RECT  3.455 2.220 3.715 2.730 ;
        RECT  2.995 2.310 3.455 2.730 ;
        RECT  2.735 2.220 2.995 2.730 ;
        RECT  1.320 2.310 2.735 2.730 ;
        RECT  1.060 2.220 1.320 2.730 ;
        RECT  0.255 2.310 1.060 2.730 ;
        RECT  0.085 1.890 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.550 0.780 6.670 1.445 ;
        RECT  6.395 0.780 6.550 0.900 ;
        RECT  6.265 1.325 6.550 1.445 ;
        RECT  6.120 1.085 6.430 1.205 ;
        RECT  6.225 0.730 6.395 0.900 ;
        RECT  6.095 1.325 6.265 1.750 ;
        RECT  6.000 0.975 6.120 1.205 ;
        RECT  5.850 1.325 6.095 1.445 ;
        RECT  5.365 0.975 6.000 1.095 ;
        RECT  5.590 1.275 5.850 1.445 ;
        RECT  5.270 0.330 5.530 0.500 ;
        RECT  5.195 0.625 5.365 1.780 ;
        RECT  5.075 0.380 5.270 0.500 ;
        RECT  5.075 1.980 5.265 2.100 ;
        RECT  4.955 0.380 5.075 2.100 ;
        RECT  4.555 0.620 4.955 0.740 ;
        RECT  2.600 1.980 4.955 2.100 ;
        RECT  4.705 1.045 4.825 1.860 ;
        RECT  3.975 1.740 4.705 1.860 ;
        RECT  4.435 0.620 4.555 1.310 ;
        RECT  4.335 1.050 4.435 1.310 ;
        RECT  4.215 1.495 4.375 1.615 ;
        RECT  4.215 0.455 4.305 0.920 ;
        RECT  4.095 0.330 4.215 1.615 ;
        RECT  3.835 0.330 4.095 0.590 ;
        RECT  3.855 0.755 3.975 1.860 ;
        RECT  3.685 0.755 3.855 0.875 ;
        RECT  2.840 1.740 3.855 1.860 ;
        RECT  3.595 1.000 3.715 1.260 ;
        RECT  3.505 1.000 3.595 1.120 ;
        RECT  3.385 0.540 3.505 1.120 ;
        RECT  2.360 0.540 3.385 0.660 ;
        RECT  2.600 0.780 3.255 0.900 ;
        RECT  2.720 1.260 2.840 1.860 ;
        RECT  2.480 0.780 2.600 2.190 ;
        RECT  2.290 2.020 2.480 2.190 ;
        RECT  2.240 0.540 2.360 1.900 ;
        RECT  2.120 2.020 2.290 2.140 ;
        RECT  2.060 0.540 2.240 0.730 ;
        RECT  2.000 0.920 2.120 2.140 ;
        RECT  1.860 0.920 2.000 1.040 ;
        RECT  1.670 0.380 1.930 0.540 ;
        RECT  1.760 1.640 1.880 2.160 ;
        RECT  0.690 1.980 1.760 2.100 ;
        RECT  0.670 0.420 1.670 0.540 ;
        RECT  0.780 0.660 1.440 0.780 ;
        RECT  0.660 0.660 0.780 1.530 ;
        RECT  0.430 1.890 0.690 2.100 ;
        RECT  0.410 0.380 0.670 0.540 ;
        RECT  0.330 0.660 0.660 0.880 ;
        RECT  0.330 1.410 0.660 1.530 ;
    END
END SDFFQXLAD
MACRO SDFFRHQX1AD
    CLASS CORE ;
    FOREIGN SDFFRHQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.900 1.140 3.930 1.400 ;
        RECT  3.810 1.015 3.900 1.400 ;
        RECT  3.710 1.015 3.810 1.375 ;
        END
        AntennaGateArea 0.05 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.080 1.390 3.200 1.660 ;
        RECT  2.580 1.540 3.080 1.660 ;
        RECT  2.460 1.280 2.580 1.660 ;
        RECT  2.225 1.280 2.460 1.400 ;
        RECT  1.985 1.175 2.225 1.400 ;
        END
        AntennaGateArea 0.103 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.760 1.175 7.880 1.635 ;
        RECT  6.970 1.175 7.760 1.295 ;
        RECT  6.710 1.080 6.970 1.375 ;
        END
        AntennaGateArea 0.105 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.410 0.640 9.450 1.565 ;
        RECT  9.290 0.640 9.410 1.895 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.675 1.160 ;
        RECT  2.265 0.900 2.350 1.050 ;
        END
        AntennaGateArea 0.084 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.025 0.530 1.375 ;
        END
        AntennaGateArea 0.114 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.090 -0.210 9.520 0.210 ;
        RECT  8.830 -0.210 9.090 0.310 ;
        RECT  8.440 -0.210 8.830 0.210 ;
        RECT  8.180 -0.210 8.440 0.310 ;
        RECT  6.760 -0.210 8.180 0.210 ;
        RECT  6.500 -0.210 6.760 0.300 ;
        RECT  5.760 -0.210 6.500 0.210 ;
        RECT  5.500 -0.210 5.760 0.300 ;
        RECT  4.415 -0.210 5.500 0.210 ;
        RECT  4.155 -0.210 4.415 0.300 ;
        RECT  2.660 -0.210 4.155 0.210 ;
        RECT  2.400 -0.210 2.660 0.300 ;
        RECT  1.425 -0.210 2.400 0.210 ;
        RECT  1.165 -0.210 1.425 0.310 ;
        RECT  0.690 -0.210 1.165 0.210 ;
        RECT  0.430 -0.210 0.690 0.310 ;
        RECT  0.000 -0.210 0.430 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.100 2.310 9.520 2.730 ;
        RECT  8.840 1.995 9.100 2.730 ;
        RECT  8.130 2.310 8.840 2.730 ;
        RECT  8.100 2.210 8.130 2.730 ;
        RECT  7.835 2.185 8.100 2.730 ;
        RECT  6.875 2.310 7.835 2.730 ;
        RECT  6.615 2.210 6.875 2.730 ;
        RECT  6.260 2.310 6.615 2.730 ;
        RECT  6.000 2.210 6.260 2.730 ;
        RECT  5.290 2.310 6.000 2.730 ;
        RECT  5.030 2.220 5.290 2.730 ;
        RECT  4.450 2.310 5.030 2.730 ;
        RECT  4.190 2.210 4.450 2.730 ;
        RECT  1.820 2.310 4.190 2.730 ;
        RECT  1.700 2.150 1.820 2.730 ;
        RECT  0.520 2.310 1.700 2.730 ;
        RECT  0.380 1.880 0.520 2.730 ;
        RECT  0.000 2.310 0.380 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.520 2.520 ;
        LAYER M1 ;
        RECT  8.930 0.520 9.050 1.875 ;
        RECT  7.955 0.520 8.930 0.640 ;
        RECT  7.480 1.755 8.930 1.875 ;
        RECT  8.740 0.760 8.810 0.880 ;
        RECT  8.620 0.760 8.740 1.590 ;
        RECT  8.550 0.760 8.620 1.070 ;
        RECT  8.360 0.950 8.550 1.070 ;
        RECT  8.350 1.330 8.470 1.590 ;
        RECT  8.240 0.950 8.360 1.210 ;
        RECT  8.120 1.330 8.350 1.450 ;
        RECT  8.000 0.935 8.120 1.450 ;
        RECT  7.210 0.935 8.000 1.055 ;
        RECT  7.835 0.520 7.955 0.815 ;
        RECT  7.450 0.695 7.835 0.815 ;
        RECT  7.330 0.555 7.450 0.815 ;
        RECT  7.240 1.440 7.380 1.560 ;
        RECT  7.210 0.330 7.260 0.450 ;
        RECT  7.120 1.440 7.240 1.720 ;
        RECT  7.090 0.330 7.210 1.055 ;
        RECT  6.590 1.600 7.120 1.720 ;
        RECT  7.000 1.930 7.120 2.190 ;
        RECT  7.000 0.330 7.090 0.540 ;
        RECT  5.270 0.420 7.000 0.540 ;
        RECT  5.750 1.970 7.000 2.090 ;
        RECT  6.800 0.680 6.970 0.850 ;
        RECT  6.590 0.680 6.800 0.800 ;
        RECT  6.470 0.680 6.590 1.845 ;
        RECT  5.860 0.680 6.470 0.800 ;
        RECT  5.350 1.220 6.470 1.340 ;
        RECT  6.385 1.600 6.470 1.845 ;
        RECT  5.220 0.980 6.200 1.100 ;
        RECT  5.490 1.970 5.750 2.180 ;
        RECT  5.370 1.650 5.630 1.830 ;
        RECT  4.410 1.970 5.490 2.090 ;
        RECT  5.220 1.650 5.370 1.770 ;
        RECT  5.010 0.350 5.270 0.540 ;
        RECT  5.095 0.730 5.220 1.770 ;
        RECT  4.860 0.730 5.095 0.850 ;
        RECT  4.680 1.650 5.095 1.770 ;
        RECT  4.005 0.420 5.010 0.540 ;
        RECT  4.730 1.150 4.830 1.410 ;
        RECT  4.610 0.660 4.730 1.410 ;
        RECT  4.560 1.590 4.680 1.850 ;
        RECT  4.170 0.660 4.610 0.780 ;
        RECT  4.410 1.080 4.450 1.340 ;
        RECT  4.290 1.080 4.410 2.090 ;
        RECT  4.060 1.970 4.290 2.090 ;
        RECT  4.050 0.660 4.170 1.850 ;
        RECT  3.940 1.970 4.060 2.140 ;
        RECT  3.485 0.660 4.050 0.780 ;
        RECT  3.820 1.730 4.050 1.850 ;
        RECT  3.885 0.380 4.005 0.540 ;
        RECT  2.060 2.020 3.940 2.140 ;
        RECT  3.215 0.380 3.885 0.500 ;
        RECT  3.560 1.730 3.820 1.900 ;
        RECT  3.440 1.480 3.635 1.600 ;
        RECT  3.320 0.940 3.440 1.900 ;
        RECT  3.170 0.940 3.320 1.060 ;
        RECT  2.300 1.780 3.320 1.900 ;
        RECT  3.005 0.660 3.310 0.780 ;
        RECT  3.095 0.380 3.215 0.540 ;
        RECT  1.870 0.420 3.095 0.540 ;
        RECT  2.960 0.660 3.005 1.225 ;
        RECT  2.885 0.660 2.960 1.420 ;
        RECT  2.790 0.660 2.885 0.780 ;
        RECT  2.840 1.105 2.885 1.420 ;
        RECT  2.700 1.300 2.840 1.420 ;
        RECT  2.180 1.520 2.300 1.900 ;
        RECT  2.140 0.660 2.280 0.780 ;
        RECT  1.865 1.520 2.180 1.640 ;
        RECT  2.020 0.660 2.140 1.055 ;
        RECT  1.940 1.820 2.060 2.140 ;
        RECT  1.865 0.935 2.020 1.055 ;
        RECT  0.770 1.820 1.940 1.990 ;
        RECT  1.750 0.420 1.870 0.815 ;
        RECT  1.745 0.935 1.865 1.640 ;
        RECT  1.625 0.695 1.750 0.815 ;
        RECT  1.505 0.695 1.625 1.635 ;
        RECT  1.010 1.465 1.505 1.635 ;
        RECT  1.265 0.495 1.385 1.285 ;
        RECT  0.375 0.495 1.265 0.615 ;
        RECT  0.890 1.135 1.010 1.635 ;
        RECT  0.770 0.735 0.935 0.905 ;
        RECT  0.650 0.735 0.770 1.990 ;
        RECT  0.265 0.495 0.375 0.855 ;
        RECT  0.255 0.495 0.265 0.905 ;
        RECT  0.210 1.495 0.265 1.665 ;
        RECT  0.210 0.735 0.255 0.905 ;
        RECT  0.090 0.735 0.210 1.665 ;
    END
END SDFFRHQX1AD
MACRO SDFFRHQX2AD
    CLASS CORE ;
    FOREIGN SDFFRHQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.900 1.140 3.930 1.400 ;
        RECT  3.810 1.015 3.900 1.400 ;
        RECT  3.710 1.015 3.810 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.080 1.390 3.200 1.660 ;
        RECT  2.580 1.540 3.080 1.660 ;
        RECT  2.460 1.280 2.580 1.660 ;
        RECT  2.225 1.280 2.460 1.400 ;
        RECT  1.985 1.175 2.225 1.400 ;
        END
        AntennaGateArea 0.118 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.760 1.175 7.880 1.635 ;
        RECT  7.010 1.175 7.760 1.295 ;
        RECT  6.790 1.000 7.010 1.375 ;
        END
        AntennaGateArea 0.141 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.290 0.385 9.450 2.020 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.350 0.900 2.675 1.160 ;
        RECT  2.265 0.900 2.350 1.050 ;
        END
        AntennaGateArea 0.132 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.050 0.530 1.655 ;
        END
        AntennaGateArea 0.119 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.050 -0.210 9.520 0.210 ;
        RECT  8.790 -0.210 9.050 0.310 ;
        RECT  8.480 -0.210 8.790 0.210 ;
        RECT  8.220 -0.210 8.480 0.310 ;
        RECT  6.750 -0.210 8.220 0.210 ;
        RECT  6.490 -0.210 6.750 0.260 ;
        RECT  5.760 -0.210 6.490 0.210 ;
        RECT  5.500 -0.210 5.760 0.260 ;
        RECT  4.415 -0.210 5.500 0.210 ;
        RECT  4.155 -0.210 4.415 0.260 ;
        RECT  2.810 -0.210 4.155 0.210 ;
        RECT  2.550 -0.210 2.810 0.300 ;
        RECT  1.420 -0.210 2.550 0.210 ;
        RECT  1.160 -0.210 1.420 0.310 ;
        RECT  0.680 -0.210 1.160 0.210 ;
        RECT  0.420 -0.210 0.680 0.310 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.100 2.310 9.520 2.730 ;
        RECT  8.840 1.995 9.100 2.730 ;
        RECT  8.130 2.310 8.840 2.730 ;
        RECT  8.100 2.210 8.130 2.730 ;
        RECT  7.835 2.185 8.100 2.730 ;
        RECT  6.830 2.310 7.835 2.730 ;
        RECT  6.660 2.265 6.830 2.730 ;
        RECT  6.200 2.310 6.660 2.730 ;
        RECT  5.940 2.220 6.200 2.730 ;
        RECT  5.380 2.310 5.940 2.730 ;
        RECT  5.120 2.220 5.380 2.730 ;
        RECT  4.450 2.310 5.120 2.730 ;
        RECT  4.190 2.210 4.450 2.730 ;
        RECT  1.820 2.310 4.190 2.730 ;
        RECT  1.700 2.150 1.820 2.730 ;
        RECT  0.520 2.310 1.700 2.730 ;
        RECT  0.380 1.900 0.520 2.730 ;
        RECT  0.000 2.310 0.380 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.520 2.520 ;
        LAYER M1 ;
        RECT  8.930 0.520 9.050 1.875 ;
        RECT  7.490 0.520 8.930 0.640 ;
        RECT  7.480 1.755 8.930 1.875 ;
        RECT  8.740 0.760 8.810 0.880 ;
        RECT  8.620 0.760 8.740 1.590 ;
        RECT  8.550 0.760 8.620 1.140 ;
        RECT  8.360 1.020 8.550 1.140 ;
        RECT  8.350 1.370 8.470 1.630 ;
        RECT  8.240 0.950 8.360 1.210 ;
        RECT  8.120 1.370 8.350 1.490 ;
        RECT  8.000 0.935 8.120 1.490 ;
        RECT  7.250 0.935 8.000 1.055 ;
        RECT  7.370 0.520 7.490 0.780 ;
        RECT  7.240 1.440 7.380 1.560 ;
        RECT  7.130 0.380 7.250 1.055 ;
        RECT  7.120 1.440 7.240 1.720 ;
        RECT  5.300 0.380 7.130 0.500 ;
        RECT  6.600 1.600 7.120 1.720 ;
        RECT  7.000 1.930 7.120 2.190 ;
        RECT  6.830 0.650 7.000 0.820 ;
        RECT  5.750 1.970 7.000 2.090 ;
        RECT  6.600 0.700 6.830 0.820 ;
        RECT  6.555 0.700 6.600 1.820 ;
        RECT  6.480 0.700 6.555 1.845 ;
        RECT  5.875 0.700 6.480 0.820 ;
        RECT  6.385 1.600 6.480 1.845 ;
        RECT  5.220 1.260 6.360 1.380 ;
        RECT  5.755 0.700 5.875 1.140 ;
        RECT  5.380 1.020 5.755 1.140 ;
        RECT  5.490 1.910 5.750 2.090 ;
        RECT  5.220 1.560 5.630 1.680 ;
        RECT  4.410 1.970 5.490 2.090 ;
        RECT  5.040 0.345 5.300 0.500 ;
        RECT  5.095 0.715 5.220 1.680 ;
        RECT  4.860 0.715 5.095 0.835 ;
        RECT  4.680 1.560 5.095 1.680 ;
        RECT  3.215 0.380 5.040 0.500 ;
        RECT  4.730 0.955 4.830 1.215 ;
        RECT  4.610 0.660 4.730 1.215 ;
        RECT  4.560 1.400 4.680 1.680 ;
        RECT  4.170 0.660 4.610 0.780 ;
        RECT  4.410 0.995 4.450 1.255 ;
        RECT  4.290 0.995 4.410 2.090 ;
        RECT  4.060 1.970 4.290 2.090 ;
        RECT  4.050 0.660 4.170 1.850 ;
        RECT  3.940 1.970 4.060 2.140 ;
        RECT  3.485 0.660 4.050 0.780 ;
        RECT  3.820 1.730 4.050 1.850 ;
        RECT  2.060 2.020 3.940 2.140 ;
        RECT  3.560 1.730 3.820 1.900 ;
        RECT  3.440 1.480 3.635 1.600 ;
        RECT  3.320 0.940 3.440 1.900 ;
        RECT  3.170 0.940 3.320 1.060 ;
        RECT  2.300 1.780 3.320 1.900 ;
        RECT  3.005 0.660 3.310 0.780 ;
        RECT  3.095 0.380 3.215 0.540 ;
        RECT  1.870 0.420 3.095 0.540 ;
        RECT  2.960 0.660 3.005 1.225 ;
        RECT  2.885 0.660 2.960 1.420 ;
        RECT  2.840 1.105 2.885 1.420 ;
        RECT  2.700 1.300 2.840 1.420 ;
        RECT  2.180 1.520 2.300 1.900 ;
        RECT  2.140 0.660 2.295 0.780 ;
        RECT  1.865 1.520 2.180 1.640 ;
        RECT  2.020 0.660 2.140 1.055 ;
        RECT  1.940 1.820 2.060 2.140 ;
        RECT  1.865 0.935 2.020 1.055 ;
        RECT  0.770 1.820 1.940 1.990 ;
        RECT  1.750 0.420 1.870 0.815 ;
        RECT  1.745 0.935 1.865 1.640 ;
        RECT  1.625 0.695 1.750 0.815 ;
        RECT  1.505 0.695 1.625 1.635 ;
        RECT  1.010 1.465 1.505 1.635 ;
        RECT  1.265 0.495 1.385 1.285 ;
        RECT  0.230 0.495 1.265 0.615 ;
        RECT  0.890 1.135 1.010 1.635 ;
        RECT  0.770 0.735 0.935 0.905 ;
        RECT  0.650 0.735 0.770 1.990 ;
        RECT  0.110 0.495 0.230 1.715 ;
    END
END SDFFRHQX2AD
MACRO SDFFRHQX4AD
    CLASS CORE ;
    FOREIGN SDFFRHQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.890 1.190 4.130 1.655 ;
        RECT  3.835 1.190 3.890 1.380 ;
        END
        AntennaGateArea 0.075 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.335 1.200 3.475 1.320 ;
        RECT  3.215 1.200 3.335 1.660 ;
        RECT  1.905 1.540 3.215 1.660 ;
        RECT  1.785 1.120 1.905 1.660 ;
        RECT  1.560 1.120 1.785 1.380 ;
        END
        AntennaGateArea 0.166 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.845 1.330 9.290 1.450 ;
        RECT  8.725 1.220 8.845 1.450 ;
        RECT  7.815 1.220 8.725 1.360 ;
        RECT  7.585 1.100 7.815 1.360 ;
        END
        AntennaGateArea 0.242 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.755 1.005 10.850 1.515 ;
        RECT  10.585 0.405 10.755 2.170 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.655 0.910 2.775 1.170 ;
        RECT  2.265 0.910 2.655 1.100 ;
        END
        AntennaGateArea 0.162 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.540 1.375 ;
        END
        AntennaGateArea 0.193 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.115 -0.210 11.200 0.210 ;
        RECT  10.945 -0.210 11.115 0.835 ;
        RECT  10.325 -0.210 10.945 0.210 ;
        RECT  10.155 -0.210 10.325 0.350 ;
        RECT  9.715 -0.210 10.155 0.210 ;
        RECT  9.545 -0.210 9.715 0.350 ;
        RECT  7.725 -0.210 9.545 0.210 ;
        RECT  7.555 -0.210 7.725 0.495 ;
        RECT  6.305 -0.210 7.555 0.210 ;
        RECT  6.045 -0.210 6.305 0.300 ;
        RECT  5.100 -0.210 6.045 0.210 ;
        RECT  4.840 -0.210 5.100 0.300 ;
        RECT  4.180 -0.210 4.840 0.210 ;
        RECT  3.920 -0.210 4.180 0.300 ;
        RECT  2.725 -0.210 3.920 0.210 ;
        RECT  2.465 -0.210 2.725 0.280 ;
        RECT  1.235 -0.210 2.465 0.210 ;
        RECT  1.065 -0.210 1.235 0.260 ;
        RECT  0.645 -0.210 1.065 0.210 ;
        RECT  0.475 -0.210 0.645 0.315 ;
        RECT  0.000 -0.210 0.475 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.115 2.310 11.200 2.730 ;
        RECT  10.945 1.730 11.115 2.730 ;
        RECT  10.385 2.310 10.945 2.730 ;
        RECT  10.215 2.020 10.385 2.730 ;
        RECT  9.385 2.310 10.215 2.730 ;
        RECT  9.215 2.010 9.385 2.730 ;
        RECT  7.595 2.310 9.215 2.730 ;
        RECT  7.425 2.210 7.595 2.730 ;
        RECT  6.880 2.310 7.425 2.730 ;
        RECT  6.620 2.210 6.880 2.730 ;
        RECT  5.590 2.310 6.620 2.730 ;
        RECT  5.330 2.210 5.590 2.730 ;
        RECT  4.590 2.310 5.330 2.730 ;
        RECT  4.330 2.260 4.590 2.730 ;
        RECT  2.665 2.310 4.330 2.730 ;
        RECT  2.405 2.260 2.665 2.730 ;
        RECT  1.955 2.310 2.405 2.730 ;
        RECT  1.695 2.260 1.955 2.730 ;
        RECT  0.585 2.310 1.695 2.730 ;
        RECT  0.415 2.030 0.585 2.730 ;
        RECT  0.000 2.310 0.415 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.200 2.520 ;
        LAYER M1 ;
        RECT  10.295 0.470 10.415 1.890 ;
        RECT  9.180 0.470 10.295 0.590 ;
        RECT  8.030 1.770 10.295 1.890 ;
        RECT  10.055 0.760 10.175 1.520 ;
        RECT  9.840 0.760 10.055 0.880 ;
        RECT  9.580 1.400 10.055 1.520 ;
        RECT  9.770 1.020 9.890 1.280 ;
        RECT  9.575 1.020 9.770 1.140 ;
        RECT  9.460 1.260 9.580 1.520 ;
        RECT  9.455 0.710 9.575 1.140 ;
        RECT  8.910 0.710 9.455 0.830 ;
        RECT  9.060 0.380 9.180 0.590 ;
        RECT  8.950 0.380 9.060 0.500 ;
        RECT  8.690 0.330 8.950 0.500 ;
        RECT  8.790 0.620 8.910 0.830 ;
        RECT  8.600 2.010 8.860 2.190 ;
        RECT  7.395 0.620 8.790 0.740 ;
        RECT  7.930 0.380 8.690 0.500 ;
        RECT  8.435 1.480 8.605 1.650 ;
        RECT  7.885 2.010 8.600 2.130 ;
        RECT  7.465 0.860 8.570 0.980 ;
        RECT  7.860 1.480 8.435 1.600 ;
        RECT  7.765 1.970 7.885 2.130 ;
        RECT  7.740 1.480 7.860 1.765 ;
        RECT  6.410 1.970 7.765 2.090 ;
        RECT  7.465 1.645 7.740 1.765 ;
        RECT  7.345 0.860 7.465 1.765 ;
        RECT  7.275 0.420 7.395 0.740 ;
        RECT  7.100 0.860 7.345 0.980 ;
        RECT  6.710 1.645 7.345 1.765 ;
        RECT  5.920 0.420 7.275 0.540 ;
        RECT  6.310 1.125 7.140 1.245 ;
        RECT  6.840 0.700 7.100 0.980 ;
        RECT  6.590 1.365 6.710 1.765 ;
        RECT  6.450 1.365 6.590 1.485 ;
        RECT  6.150 1.970 6.410 2.190 ;
        RECT  6.190 0.680 6.310 1.845 ;
        RECT  5.620 0.680 6.190 0.800 ;
        RECT  4.890 1.725 6.190 1.845 ;
        RECT  4.610 1.970 6.150 2.090 ;
        RECT  5.910 1.340 6.070 1.460 ;
        RECT  5.660 0.350 5.920 0.540 ;
        RECT  5.780 1.110 5.910 1.460 ;
        RECT  5.070 1.110 5.780 1.230 ;
        RECT  3.750 0.420 5.660 0.540 ;
        RECT  5.500 0.660 5.620 0.800 ;
        RECT  4.180 0.660 5.500 0.780 ;
        RECT  4.950 0.925 5.070 1.230 ;
        RECT  4.370 0.925 4.950 1.045 ;
        RECT  4.770 1.585 4.890 1.845 ;
        RECT  4.610 1.255 4.795 1.375 ;
        RECT  4.490 1.255 4.610 2.140 ;
        RECT  1.170 2.020 4.490 2.140 ;
        RECT  4.250 0.925 4.370 1.900 ;
        RECT  3.990 0.925 4.250 1.045 ;
        RECT  3.695 1.780 4.250 1.900 ;
        RECT  3.865 0.660 3.990 1.045 ;
        RECT  3.550 0.660 3.865 0.780 ;
        RECT  3.715 1.500 3.770 1.620 ;
        RECT  3.630 0.400 3.750 0.540 ;
        RECT  3.595 0.960 3.715 1.620 ;
        RECT  2.585 0.400 3.630 0.520 ;
        RECT  3.410 0.960 3.595 1.080 ;
        RECT  3.575 1.500 3.595 1.620 ;
        RECT  3.455 1.500 3.575 1.900 ;
        RECT  3.290 0.640 3.550 0.780 ;
        RECT  1.665 1.780 3.455 1.900 ;
        RECT  3.150 0.900 3.410 1.080 ;
        RECT  3.015 0.640 3.170 0.760 ;
        RECT  3.015 1.300 3.095 1.420 ;
        RECT  2.895 0.640 3.015 1.420 ;
        RECT  2.835 1.300 2.895 1.420 ;
        RECT  2.465 0.400 2.585 0.740 ;
        RECT  2.145 0.620 2.465 0.740 ;
        RECT  2.145 1.300 2.395 1.420 ;
        RECT  2.025 0.620 2.145 1.420 ;
        RECT  0.945 0.380 2.040 0.500 ;
        RECT  1.175 0.620 2.025 0.740 ;
        RECT  1.440 0.860 1.700 0.980 ;
        RECT  1.545 1.555 1.665 1.900 ;
        RECT  1.440 1.555 1.545 1.675 ;
        RECT  1.320 0.860 1.440 1.675 ;
        RECT  1.055 0.620 1.175 1.260 ;
        RECT  1.050 1.460 1.170 2.140 ;
        RECT  0.900 1.140 1.055 1.260 ;
        RECT  0.780 1.460 1.050 1.580 ;
        RECT  0.825 0.380 0.945 0.555 ;
        RECT  0.800 0.675 0.920 0.935 ;
        RECT  0.230 0.435 0.825 0.555 ;
        RECT  0.780 0.810 0.800 0.935 ;
        RECT  0.660 0.810 0.780 1.580 ;
        RECT  0.110 0.435 0.230 1.730 ;
    END
END SDFFRHQX4AD
MACRO SDFFRHQX8AD
    CLASS CORE ;
    FOREIGN SDFFRHQX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.200 1.165 4.555 1.380 ;
        END
        AntennaGateArea 0.118 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.675 1.150 3.795 1.660 ;
        RECT  2.365 1.540 3.675 1.660 ;
        RECT  2.245 1.120 2.365 1.660 ;
        RECT  2.020 1.120 2.245 1.375 ;
        END
        AntennaGateArea 0.188 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.490 1.220 9.750 1.390 ;
        RECT  8.375 1.220 9.490 1.360 ;
        RECT  7.980 1.100 8.375 1.360 ;
        END
        AntennaGateArea 0.293 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.705 0.365 11.875 2.170 ;
        RECT  11.155 1.005 11.705 1.515 ;
        RECT  10.985 0.365 11.155 2.170 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.155 0.910 3.275 1.170 ;
        RECT  2.825 0.910 3.155 1.100 ;
        END
        AntennaGateArea 0.158 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.540 1.375 ;
        END
        AntennaGateArea 0.353 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.235 -0.210 12.320 0.210 ;
        RECT  12.065 -0.210 12.235 0.795 ;
        RECT  11.515 -0.210 12.065 0.210 ;
        RECT  11.345 -0.210 11.515 0.795 ;
        RECT  10.725 -0.210 11.345 0.210 ;
        RECT  10.555 -0.210 10.725 0.350 ;
        RECT  10.235 -0.210 10.555 0.210 ;
        RECT  10.065 -0.210 10.235 0.350 ;
        RECT  8.185 -0.210 10.065 0.210 ;
        RECT  8.015 -0.210 8.185 0.500 ;
        RECT  6.765 -0.210 8.015 0.210 ;
        RECT  6.505 -0.210 6.765 0.300 ;
        RECT  5.560 -0.210 6.505 0.210 ;
        RECT  5.300 -0.210 5.560 0.300 ;
        RECT  4.645 -0.210 5.300 0.210 ;
        RECT  4.385 -0.210 4.645 0.300 ;
        RECT  3.275 -0.210 4.385 0.210 ;
        RECT  3.015 -0.210 3.275 0.260 ;
        RECT  2.440 -0.210 3.015 0.210 ;
        RECT  2.440 0.330 2.490 0.500 ;
        RECT  2.320 -0.210 2.440 0.500 ;
        RECT  1.645 -0.210 2.320 0.210 ;
        RECT  1.475 -0.210 1.645 0.260 ;
        RECT  0.660 -0.210 1.475 0.210 ;
        RECT  0.400 -0.210 0.660 0.400 ;
        RECT  0.000 -0.210 0.400 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.210 2.310 12.320 2.730 ;
        RECT  12.090 1.435 12.210 2.730 ;
        RECT  11.515 2.310 12.090 2.730 ;
        RECT  11.345 1.730 11.515 2.730 ;
        RECT  10.770 2.310 11.345 2.730 ;
        RECT  10.510 2.210 10.770 2.730 ;
        RECT  9.880 2.310 10.510 2.730 ;
        RECT  9.620 2.120 9.880 2.730 ;
        RECT  8.055 2.310 9.620 2.730 ;
        RECT  7.885 2.265 8.055 2.730 ;
        RECT  7.340 2.310 7.885 2.730 ;
        RECT  7.080 2.210 7.340 2.730 ;
        RECT  6.050 2.310 7.080 2.730 ;
        RECT  5.790 2.210 6.050 2.730 ;
        RECT  5.095 2.310 5.790 2.730 ;
        RECT  4.835 2.260 5.095 2.730 ;
        RECT  3.125 2.310 4.835 2.730 ;
        RECT  2.865 2.290 3.125 2.730 ;
        RECT  2.410 2.310 2.865 2.730 ;
        RECT  2.240 2.260 2.410 2.730 ;
        RECT  1.905 2.310 2.240 2.730 ;
        RECT  1.735 2.260 1.905 2.730 ;
        RECT  0.615 2.310 1.735 2.730 ;
        RECT  0.445 1.855 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 12.320 2.520 ;
        LAYER M1 ;
        RECT  10.745 0.470 10.865 2.000 ;
        RECT  9.705 0.470 10.745 0.590 ;
        RECT  9.615 1.880 10.745 2.000 ;
        RECT  10.470 0.760 10.590 1.520 ;
        RECT  10.270 0.760 10.470 0.880 ;
        RECT  10.110 1.400 10.470 1.520 ;
        RECT  10.230 1.020 10.350 1.280 ;
        RECT  10.035 1.020 10.230 1.140 ;
        RECT  9.990 1.400 10.110 1.760 ;
        RECT  9.915 0.710 10.035 1.140 ;
        RECT  9.870 1.500 9.990 1.760 ;
        RECT  9.370 0.710 9.915 0.830 ;
        RECT  9.585 0.380 9.705 0.590 ;
        RECT  9.495 1.770 9.615 2.000 ;
        RECT  9.390 0.380 9.585 0.500 ;
        RECT  8.450 1.770 9.495 1.890 ;
        RECT  9.130 0.330 9.390 0.500 ;
        RECT  9.250 0.620 9.370 0.830 ;
        RECT  9.060 2.010 9.320 2.190 ;
        RECT  7.855 0.620 9.250 0.740 ;
        RECT  8.565 0.380 9.130 0.500 ;
        RECT  8.895 1.480 9.065 1.650 ;
        RECT  8.345 2.010 9.060 2.130 ;
        RECT  7.840 0.860 9.005 0.980 ;
        RECT  8.320 1.480 8.895 1.600 ;
        RECT  8.395 0.330 8.565 0.500 ;
        RECT  8.225 1.970 8.345 2.130 ;
        RECT  8.200 1.480 8.320 1.765 ;
        RECT  6.870 1.970 8.225 2.090 ;
        RECT  7.840 1.645 8.200 1.765 ;
        RECT  7.735 0.420 7.855 0.740 ;
        RECT  7.720 0.860 7.840 1.765 ;
        RECT  6.380 0.420 7.735 0.540 ;
        RECT  7.560 0.860 7.720 0.980 ;
        RECT  7.170 1.645 7.720 1.765 ;
        RECT  6.770 1.125 7.600 1.245 ;
        RECT  7.300 0.700 7.560 0.980 ;
        RECT  7.050 1.365 7.170 1.765 ;
        RECT  6.910 1.365 7.050 1.485 ;
        RECT  6.610 1.970 6.870 2.190 ;
        RECT  6.650 0.680 6.770 1.845 ;
        RECT  6.080 0.680 6.650 0.800 ;
        RECT  5.350 1.725 6.650 1.845 ;
        RECT  5.110 1.970 6.610 2.090 ;
        RECT  6.370 1.320 6.530 1.440 ;
        RECT  6.120 0.350 6.380 0.540 ;
        RECT  6.240 1.110 6.370 1.440 ;
        RECT  5.530 1.110 6.240 1.230 ;
        RECT  4.210 0.420 6.120 0.540 ;
        RECT  5.960 0.660 6.080 0.800 ;
        RECT  4.640 0.660 5.960 0.780 ;
        RECT  5.410 0.925 5.530 1.230 ;
        RECT  4.870 0.925 5.410 1.045 ;
        RECT  5.230 1.585 5.350 1.845 ;
        RECT  5.110 1.255 5.255 1.375 ;
        RECT  4.990 1.255 5.110 2.140 ;
        RECT  1.855 2.020 4.990 2.140 ;
        RECT  4.750 0.925 4.870 1.900 ;
        RECT  4.450 0.925 4.750 1.045 ;
        RECT  4.155 1.780 4.750 1.900 ;
        RECT  4.325 0.670 4.450 1.045 ;
        RECT  3.970 0.670 4.325 0.790 ;
        RECT  4.090 0.380 4.210 0.540 ;
        RECT  4.035 1.520 4.175 1.640 ;
        RECT  3.235 0.380 4.090 0.500 ;
        RECT  3.915 0.910 4.035 1.900 ;
        RECT  3.800 0.620 3.970 0.790 ;
        RECT  3.635 0.910 3.915 1.030 ;
        RECT  2.095 1.780 3.915 1.900 ;
        RECT  3.515 0.620 3.610 0.790 ;
        RECT  3.515 1.300 3.555 1.420 ;
        RECT  3.395 0.620 3.515 1.420 ;
        RECT  3.295 1.300 3.395 1.420 ;
        RECT  3.115 0.380 3.235 0.740 ;
        RECT  2.605 0.620 3.115 0.740 ;
        RECT  2.605 1.300 2.855 1.420 ;
        RECT  2.485 0.620 2.605 1.420 ;
        RECT  1.300 0.620 2.485 0.740 ;
        RECT  1.940 0.330 2.200 0.500 ;
        RECT  1.900 0.860 2.160 0.980 ;
        RECT  1.975 1.495 2.095 1.900 ;
        RECT  1.900 1.495 1.975 1.615 ;
        RECT  0.900 0.380 1.940 0.500 ;
        RECT  1.780 0.860 1.900 1.615 ;
        RECT  1.735 1.865 1.855 2.140 ;
        RECT  1.200 1.865 1.735 1.985 ;
        RECT  1.180 0.620 1.300 1.400 ;
        RECT  1.080 1.620 1.200 2.140 ;
        RECT  1.040 1.280 1.180 1.400 ;
        RECT  0.780 1.620 1.080 1.740 ;
        RECT  0.780 0.760 1.040 0.880 ;
        RECT  0.780 0.380 0.900 0.640 ;
        RECT  0.230 0.520 0.780 0.640 ;
        RECT  0.660 0.760 0.780 1.740 ;
        RECT  0.110 0.330 0.230 1.965 ;
    END
END SDFFRHQX8AD
MACRO SDFFRQX1AD
    CLASS CORE ;
    FOREIGN SDFFRQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.865 1.630 1.530 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.705 0.430 1.935 ;
        END
        AntennaGateArea 0.106 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.460 0.990 6.610 1.250 ;
        RECT  6.160 0.990 6.460 1.110 ;
        RECT  6.040 0.415 6.160 1.110 ;
        RECT  5.450 0.415 6.040 0.535 ;
        RECT  5.330 0.415 5.450 0.685 ;
        RECT  4.870 0.565 5.330 0.685 ;
        RECT  4.810 0.565 4.870 0.840 ;
        RECT  4.690 0.380 4.810 0.840 ;
        RECT  3.170 0.380 4.690 0.500 ;
        RECT  3.050 0.380 3.170 0.540 ;
        RECT  2.450 0.420 3.050 0.540 ;
        RECT  2.330 0.420 2.450 0.935 ;
        RECT  2.190 0.815 2.330 0.935 ;
        RECT  2.150 0.815 2.190 1.095 ;
        RECT  2.030 0.815 2.150 1.390 ;
        RECT  2.025 1.270 2.030 1.390 ;
        RECT  1.855 1.270 2.025 1.560 ;
        END
        AntennaGateArea 0.124 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.730 0.330 7.770 1.555 ;
        RECT  7.610 0.330 7.730 1.945 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.110 0.870 1.450 ;
        END
        AntennaGateArea 0.065 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.055 2.575 1.375 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.440 -0.210 7.840 0.210 ;
        RECT  7.180 -0.210 7.440 0.470 ;
        RECT  6.455 -0.210 7.180 0.210 ;
        RECT  6.285 -0.210 6.455 0.840 ;
        RECT  5.210 -0.210 6.285 0.210 ;
        RECT  4.950 -0.210 5.210 0.445 ;
        RECT  2.940 -0.210 4.950 0.210 ;
        RECT  2.420 -0.210 2.940 0.300 ;
        RECT  0.230 -0.210 2.420 0.210 ;
        RECT  0.110 -0.210 0.230 0.940 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.420 2.310 7.840 2.730 ;
        RECT  7.250 1.425 7.420 2.730 ;
        RECT  6.575 2.310 7.250 2.730 ;
        RECT  6.405 1.855 6.575 2.730 ;
        RECT  4.540 2.310 6.405 2.730 ;
        RECT  4.280 2.095 4.540 2.730 ;
        RECT  2.860 2.310 4.280 2.730 ;
        RECT  2.600 2.220 2.860 2.730 ;
        RECT  1.765 2.310 2.600 2.730 ;
        RECT  1.595 2.175 1.765 2.730 ;
        RECT  0.600 2.310 1.595 2.730 ;
        RECT  0.340 2.055 0.600 2.730 ;
        RECT  0.000 2.310 0.340 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.840 2.520 ;
        LAYER M1 ;
        RECT  7.310 0.755 7.480 1.185 ;
        RECT  7.130 0.985 7.310 1.185 ;
        RECT  7.010 0.695 7.130 1.735 ;
        RECT  6.850 0.695 7.010 0.815 ;
        RECT  6.240 1.615 7.010 1.735 ;
        RECT  6.770 0.995 6.890 1.490 ;
        RECT  5.780 1.370 6.770 1.490 ;
        RECT  6.120 1.615 6.240 2.115 ;
        RECT  5.830 2.070 5.970 2.190 ;
        RECT  5.780 0.670 5.845 0.840 ;
        RECT  5.710 1.925 5.830 2.190 ;
        RECT  5.660 0.670 5.780 1.805 ;
        RECT  5.060 1.925 5.710 2.045 ;
        RECT  5.620 1.545 5.660 1.805 ;
        RECT  5.295 0.805 5.465 1.760 ;
        RECT  5.235 1.270 5.295 1.760 ;
        RECT  4.640 1.270 5.235 1.390 ;
        RECT  4.940 1.585 5.060 2.045 ;
        RECT  4.400 1.585 4.940 1.705 ;
        RECT  4.700 1.855 4.820 2.120 ;
        RECT  4.160 1.855 4.700 1.975 ;
        RECT  4.520 1.205 4.640 1.465 ;
        RECT  4.280 0.620 4.400 1.705 ;
        RECT  3.540 0.620 4.280 0.740 ;
        RECT  4.040 0.890 4.160 2.100 ;
        RECT  1.930 1.980 4.040 2.100 ;
        RECT  3.750 0.890 3.870 1.860 ;
        RECT  3.660 0.890 3.750 1.150 ;
        RECT  1.350 1.740 3.750 1.860 ;
        RECT  3.420 0.620 3.540 1.560 ;
        RECT  3.340 0.620 3.420 0.740 ;
        RECT  2.935 1.390 3.420 1.560 ;
        RECT  3.180 0.885 3.300 1.145 ;
        RECT  2.815 1.025 3.180 1.145 ;
        RECT  2.815 0.660 2.880 0.780 ;
        RECT  2.695 0.660 2.815 1.615 ;
        RECT  2.620 0.660 2.695 0.780 ;
        RECT  2.220 1.495 2.695 1.615 ;
        RECT  1.955 0.380 2.125 0.695 ;
        RECT  0.865 0.380 1.955 0.500 ;
        RECT  1.350 0.620 1.540 0.740 ;
        RECT  1.230 0.620 1.350 1.860 ;
        RECT  1.025 1.660 1.230 1.860 ;
        RECT  0.990 0.840 1.110 1.360 ;
        RECT  0.660 0.840 0.990 0.960 ;
        RECT  0.695 0.380 0.865 0.555 ;
        RECT  0.470 0.750 0.660 0.960 ;
        RECT  0.400 0.750 0.470 1.180 ;
        RECT  0.350 0.840 0.400 1.180 ;
        RECT  0.255 1.060 0.350 1.180 ;
        RECT  0.135 1.060 0.255 1.555 ;
        RECT  0.085 1.385 0.135 1.555 ;
    END
END SDFFRQX1AD
MACRO SDFFRQX2AD
    CLASS CORE ;
    FOREIGN SDFFRQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.660 0.865 1.890 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.705 0.355 2.020 ;
        RECT  0.070 1.705 0.185 1.935 ;
        END
        AntennaGateArea 0.105 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.435 0.330 6.605 0.580 ;
        RECT  5.250 0.380 6.435 0.500 ;
        RECT  5.130 0.380 5.250 0.785 ;
        RECT  5.080 0.665 5.130 0.785 ;
        RECT  4.820 0.665 5.080 1.155 ;
        RECT  4.725 0.665 4.820 0.785 ;
        RECT  4.605 0.380 4.725 0.785 ;
        RECT  3.155 0.380 4.605 0.500 ;
        RECT  3.035 0.380 3.155 0.540 ;
        RECT  2.450 0.420 3.035 0.540 ;
        RECT  2.330 0.420 2.450 1.020 ;
        RECT  2.140 0.900 2.330 1.020 ;
        RECT  2.020 0.900 2.140 1.585 ;
        END
        AntennaGateArea 0.13 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.610 0.365 7.770 2.030 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.605 1.110 0.910 1.375 ;
        END
        AntennaGateArea 0.064 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.580 1.020 2.700 1.375 ;
        RECT  2.310 1.145 2.580 1.375 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.395 -0.210 7.840 0.210 ;
        RECT  7.225 -0.210 7.395 0.535 ;
        RECT  6.845 -0.210 7.225 0.210 ;
        RECT  6.725 -0.210 6.845 0.820 ;
        RECT  5.010 -0.210 6.725 0.210 ;
        RECT  6.270 0.700 6.725 0.820 ;
        RECT  4.890 -0.210 5.010 0.505 ;
        RECT  2.925 -0.210 4.890 0.210 ;
        RECT  2.405 -0.210 2.925 0.300 ;
        RECT  0.230 -0.210 2.405 0.210 ;
        RECT  0.110 -0.210 0.230 0.940 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.420 2.310 7.840 2.730 ;
        RECT  7.250 1.510 7.420 2.730 ;
        RECT  6.415 2.310 7.250 2.730 ;
        RECT  6.245 2.020 6.415 2.730 ;
        RECT  5.010 2.310 6.245 2.730 ;
        RECT  4.840 1.825 5.010 2.730 ;
        RECT  4.445 2.310 4.840 2.730 ;
        RECT  4.185 2.105 4.445 2.730 ;
        RECT  2.900 2.310 4.185 2.730 ;
        RECT  2.640 2.220 2.900 2.730 ;
        RECT  1.960 2.310 2.640 2.730 ;
        RECT  1.700 1.980 1.960 2.730 ;
        RECT  0.645 2.310 1.700 2.730 ;
        RECT  0.475 1.505 0.645 2.730 ;
        RECT  0.000 2.310 0.475 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.840 2.520 ;
        LAYER M1 ;
        RECT  7.130 1.020 7.470 1.280 ;
        RECT  7.010 0.630 7.130 1.735 ;
        RECT  6.965 0.630 7.010 0.890 ;
        RECT  6.310 1.615 7.010 1.735 ;
        RECT  6.860 1.235 6.890 1.495 ;
        RECT  6.740 0.990 6.860 1.495 ;
        RECT  5.875 0.990 6.740 1.110 ;
        RECT  6.190 1.235 6.310 1.735 ;
        RECT  5.815 1.925 6.075 2.190 ;
        RECT  5.755 0.675 5.875 1.760 ;
        RECT  5.250 1.925 5.815 2.045 ;
        RECT  5.705 0.675 5.755 0.845 ;
        RECT  5.705 1.590 5.755 1.760 ;
        RECT  5.370 0.630 5.490 1.805 ;
        RECT  4.605 1.335 5.370 1.455 ;
        RECT  5.130 1.585 5.250 2.045 ;
        RECT  4.485 1.585 5.130 1.705 ;
        RECT  4.595 1.865 4.715 2.125 ;
        RECT  4.240 1.865 4.595 1.985 ;
        RECT  4.365 0.620 4.485 1.705 ;
        RECT  3.600 0.620 4.365 0.740 ;
        RECT  4.120 0.860 4.240 1.985 ;
        RECT  3.910 1.865 4.120 1.985 ;
        RECT  3.860 1.730 3.910 1.985 ;
        RECT  3.840 0.860 3.880 1.120 ;
        RECT  3.740 1.730 3.860 2.100 ;
        RECT  3.720 0.860 3.840 1.610 ;
        RECT  2.080 1.980 3.740 2.100 ;
        RECT  3.595 1.490 3.720 1.610 ;
        RECT  3.480 0.620 3.600 1.370 ;
        RECT  3.475 1.490 3.595 1.860 ;
        RECT  3.270 0.660 3.480 0.780 ;
        RECT  3.220 1.250 3.480 1.370 ;
        RECT  1.530 1.740 3.475 1.860 ;
        RECT  2.955 0.945 3.295 1.115 ;
        RECT  3.100 1.250 3.220 1.605 ;
        RECT  2.835 0.660 2.955 1.615 ;
        RECT  2.600 0.660 2.835 0.780 ;
        RECT  2.360 1.495 2.835 1.615 ;
        RECT  2.100 0.610 2.150 0.780 ;
        RECT  1.980 0.380 2.100 0.780 ;
        RECT  0.895 0.380 1.980 0.500 ;
        RECT  1.530 0.635 1.580 0.755 ;
        RECT  1.410 0.635 1.530 1.860 ;
        RECT  1.320 0.635 1.410 0.755 ;
        RECT  1.105 1.665 1.410 1.860 ;
        RECT  1.150 1.155 1.290 1.275 ;
        RECT  1.030 0.840 1.150 1.275 ;
        RECT  0.615 0.840 1.030 0.960 ;
        RECT  0.725 0.380 0.895 0.555 ;
        RECT  0.480 0.725 0.615 0.960 ;
        RECT  0.445 0.725 0.480 1.180 ;
        RECT  0.360 0.840 0.445 1.180 ;
        RECT  0.255 1.060 0.360 1.180 ;
        RECT  0.135 1.060 0.255 1.555 ;
        RECT  0.085 1.385 0.135 1.555 ;
    END
END SDFFRQX2AD
MACRO SDFFRQX4AD
    CLASS CORE ;
    FOREIGN SDFFRQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.660 0.865 1.890 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.705 0.355 2.020 ;
        RECT  0.070 1.705 0.185 1.935 ;
        END
        AntennaGateArea 0.105 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.360 0.980 6.870 1.100 ;
        RECT  6.240 0.380 6.360 1.100 ;
        RECT  5.420 0.380 6.240 0.500 ;
        RECT  5.300 0.380 5.420 0.785 ;
        RECT  5.250 0.665 5.300 0.785 ;
        RECT  4.990 0.665 5.250 1.155 ;
        RECT  4.895 0.665 4.990 0.785 ;
        RECT  4.775 0.380 4.895 0.785 ;
        RECT  3.475 0.380 4.775 0.500 ;
        RECT  3.355 0.380 3.475 0.540 ;
        RECT  2.450 0.420 3.355 0.540 ;
        RECT  2.330 0.420 2.450 1.115 ;
        RECT  2.220 0.945 2.330 1.115 ;
        RECT  2.175 0.995 2.220 1.115 ;
        RECT  2.055 0.995 2.175 1.595 ;
        RECT  2.005 1.425 2.055 1.595 ;
        END
        AntennaGateArea 0.167 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.960 0.880 8.050 1.625 ;
        RECT  7.800 0.365 7.960 2.030 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.605 1.110 0.910 1.375 ;
        END
        AntennaGateArea 0.064 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.900 2.775 1.375 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.305 -0.210 8.400 0.210 ;
        RECT  8.135 -0.210 8.305 0.510 ;
        RECT  7.585 -0.210 8.135 0.210 ;
        RECT  7.415 -0.210 7.585 0.510 ;
        RECT  6.740 -0.210 7.415 0.210 ;
        RECT  6.480 -0.210 6.740 0.820 ;
        RECT  5.180 -0.210 6.480 0.210 ;
        RECT  5.060 -0.210 5.180 0.505 ;
        RECT  3.220 -0.210 5.060 0.210 ;
        RECT  2.960 -0.210 3.220 0.300 ;
        RECT  2.575 -0.210 2.960 0.210 ;
        RECT  2.315 -0.210 2.575 0.300 ;
        RECT  0.230 -0.210 2.315 0.210 ;
        RECT  0.110 -0.210 0.230 0.940 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.305 2.310 8.400 2.730 ;
        RECT  8.135 1.845 8.305 2.730 ;
        RECT  7.585 2.310 8.135 2.730 ;
        RECT  7.415 1.845 7.585 2.730 ;
        RECT  6.705 2.310 7.415 2.730 ;
        RECT  6.535 1.715 6.705 2.730 ;
        RECT  4.865 2.310 6.535 2.730 ;
        RECT  4.605 2.105 4.865 2.730 ;
        RECT  3.075 2.310 4.605 2.730 ;
        RECT  2.815 2.220 3.075 2.730 ;
        RECT  1.960 2.310 2.815 2.730 ;
        RECT  1.700 1.980 1.960 2.730 ;
        RECT  0.645 2.310 1.700 2.730 ;
        RECT  0.475 1.505 0.645 2.730 ;
        RECT  0.000 2.310 0.475 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.400 2.520 ;
        LAYER M1 ;
        RECT  7.450 1.020 7.660 1.280 ;
        RECT  7.330 0.675 7.450 1.580 ;
        RECT  7.145 0.675 7.330 0.845 ;
        RECT  7.065 1.460 7.330 1.580 ;
        RECT  7.025 1.145 7.195 1.340 ;
        RECT  6.895 1.460 7.065 2.010 ;
        RECT  6.095 1.220 7.025 1.340 ;
        RECT  6.360 1.460 6.895 1.580 ;
        RECT  5.990 1.925 6.250 2.190 ;
        RECT  5.895 0.675 6.095 1.685 ;
        RECT  5.420 1.925 5.990 2.045 ;
        RECT  5.560 0.630 5.680 1.780 ;
        RECT  4.775 1.335 5.560 1.455 ;
        RECT  5.300 1.585 5.420 2.045 ;
        RECT  4.655 1.585 5.300 1.705 ;
        RECT  5.010 1.865 5.130 2.125 ;
        RECT  4.410 1.865 5.010 1.985 ;
        RECT  4.535 0.620 4.655 1.705 ;
        RECT  3.725 0.620 4.535 0.740 ;
        RECT  4.290 0.860 4.410 1.985 ;
        RECT  4.120 1.730 4.290 1.985 ;
        RECT  4.000 1.730 4.120 2.100 ;
        RECT  4.010 0.860 4.050 1.120 ;
        RECT  3.890 0.860 4.010 1.610 ;
        RECT  2.080 1.980 4.000 2.100 ;
        RECT  3.855 1.490 3.890 1.610 ;
        RECT  3.735 1.490 3.855 1.860 ;
        RECT  1.530 1.740 3.735 1.860 ;
        RECT  3.605 0.620 3.725 1.355 ;
        RECT  3.340 0.660 3.605 0.780 ;
        RECT  3.555 1.185 3.605 1.355 ;
        RECT  3.410 1.235 3.555 1.355 ;
        RECT  3.290 1.235 3.410 1.605 ;
        RECT  3.095 0.945 3.315 1.115 ;
        RECT  2.975 0.660 3.095 1.615 ;
        RECT  2.600 0.660 2.975 0.780 ;
        RECT  2.435 1.495 2.975 1.615 ;
        RECT  2.100 0.610 2.150 0.780 ;
        RECT  1.980 0.380 2.100 0.780 ;
        RECT  0.895 0.380 1.980 0.500 ;
        RECT  1.530 0.635 1.580 0.755 ;
        RECT  1.410 0.635 1.530 1.860 ;
        RECT  1.320 0.635 1.410 0.755 ;
        RECT  1.105 1.665 1.410 1.860 ;
        RECT  1.150 1.155 1.290 1.275 ;
        RECT  1.030 0.840 1.150 1.275 ;
        RECT  0.615 0.840 1.030 0.960 ;
        RECT  0.725 0.380 0.895 0.555 ;
        RECT  0.480 0.725 0.615 0.960 ;
        RECT  0.445 0.725 0.480 1.180 ;
        RECT  0.360 0.840 0.445 1.180 ;
        RECT  0.255 1.060 0.360 1.180 ;
        RECT  0.135 1.060 0.255 1.555 ;
        RECT  0.085 1.385 0.135 1.555 ;
    END
END SDFFRQX4AD
MACRO SDFFRQXLAD
    CLASS CORE ;
    FOREIGN SDFFRQXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.865 1.630 1.530 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.705 0.430 1.935 ;
        END
        AntennaGateArea 0.106 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.460 0.990 6.610 1.250 ;
        RECT  6.160 0.990 6.460 1.110 ;
        RECT  6.040 0.415 6.160 1.110 ;
        RECT  5.450 0.415 6.040 0.535 ;
        RECT  5.330 0.415 5.450 0.685 ;
        RECT  4.870 0.565 5.330 0.685 ;
        RECT  4.810 0.565 4.870 0.840 ;
        RECT  4.690 0.380 4.810 0.840 ;
        RECT  3.170 0.380 4.690 0.500 ;
        RECT  3.050 0.380 3.170 0.540 ;
        RECT  2.450 0.420 3.050 0.540 ;
        RECT  2.330 0.420 2.450 0.935 ;
        RECT  2.190 0.815 2.330 0.935 ;
        RECT  2.150 0.815 2.190 1.095 ;
        RECT  2.030 0.815 2.150 1.390 ;
        RECT  2.025 1.270 2.030 1.390 ;
        RECT  1.855 1.270 2.025 1.560 ;
        END
        AntennaGateArea 0.124 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.610 0.330 7.770 1.710 ;
        END
        AntennaDiffArea 0.143 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.110 0.870 1.450 ;
        END
        AntennaGateArea 0.065 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.055 2.575 1.375 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.440 -0.210 7.840 0.210 ;
        RECT  7.180 -0.210 7.440 0.520 ;
        RECT  6.455 -0.210 7.180 0.210 ;
        RECT  6.285 -0.210 6.455 0.840 ;
        RECT  5.210 -0.210 6.285 0.210 ;
        RECT  4.950 -0.210 5.210 0.445 ;
        RECT  2.940 -0.210 4.950 0.210 ;
        RECT  2.420 -0.210 2.940 0.300 ;
        RECT  0.230 -0.210 2.420 0.210 ;
        RECT  0.110 -0.210 0.230 0.940 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.420 2.310 7.840 2.730 ;
        RECT  7.250 1.425 7.420 2.730 ;
        RECT  6.575 2.310 7.250 2.730 ;
        RECT  6.405 1.855 6.575 2.730 ;
        RECT  4.540 2.310 6.405 2.730 ;
        RECT  4.280 2.095 4.540 2.730 ;
        RECT  2.860 2.310 4.280 2.730 ;
        RECT  2.600 2.220 2.860 2.730 ;
        RECT  1.765 2.310 2.600 2.730 ;
        RECT  1.595 2.175 1.765 2.730 ;
        RECT  0.600 2.310 1.595 2.730 ;
        RECT  0.340 2.055 0.600 2.730 ;
        RECT  0.000 2.310 0.340 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.840 2.520 ;
        LAYER M1 ;
        RECT  7.310 0.755 7.480 1.185 ;
        RECT  7.130 0.985 7.310 1.185 ;
        RECT  7.010 0.695 7.130 1.735 ;
        RECT  6.850 0.695 7.010 0.815 ;
        RECT  6.240 1.615 7.010 1.735 ;
        RECT  6.770 0.995 6.890 1.490 ;
        RECT  5.780 1.370 6.770 1.490 ;
        RECT  6.120 1.615 6.240 2.115 ;
        RECT  5.830 2.070 5.970 2.190 ;
        RECT  5.780 0.670 5.845 0.840 ;
        RECT  5.710 1.925 5.830 2.190 ;
        RECT  5.660 0.670 5.780 1.805 ;
        RECT  5.060 1.925 5.710 2.045 ;
        RECT  5.620 1.545 5.660 1.805 ;
        RECT  5.295 0.805 5.465 1.760 ;
        RECT  5.235 1.270 5.295 1.760 ;
        RECT  4.640 1.270 5.235 1.390 ;
        RECT  4.940 1.585 5.060 2.045 ;
        RECT  4.400 1.585 4.940 1.705 ;
        RECT  4.700 1.855 4.820 2.120 ;
        RECT  4.160 1.855 4.700 1.975 ;
        RECT  4.520 1.205 4.640 1.465 ;
        RECT  4.280 0.620 4.400 1.705 ;
        RECT  3.540 0.620 4.280 0.740 ;
        RECT  4.040 0.890 4.160 2.100 ;
        RECT  1.930 1.980 4.040 2.100 ;
        RECT  3.750 0.890 3.870 1.860 ;
        RECT  3.660 0.890 3.750 1.150 ;
        RECT  1.350 1.740 3.750 1.860 ;
        RECT  3.420 0.620 3.540 1.560 ;
        RECT  3.340 0.620 3.420 0.740 ;
        RECT  2.935 1.390 3.420 1.560 ;
        RECT  3.180 0.885 3.300 1.145 ;
        RECT  2.815 1.025 3.180 1.145 ;
        RECT  2.815 0.660 2.880 0.780 ;
        RECT  2.695 0.660 2.815 1.615 ;
        RECT  2.620 0.660 2.695 0.780 ;
        RECT  2.220 1.495 2.695 1.615 ;
        RECT  1.955 0.380 2.125 0.695 ;
        RECT  0.865 0.380 1.955 0.500 ;
        RECT  1.350 0.620 1.540 0.740 ;
        RECT  1.230 0.620 1.350 1.860 ;
        RECT  1.025 1.660 1.230 1.860 ;
        RECT  0.990 0.840 1.110 1.360 ;
        RECT  0.660 0.840 0.990 0.960 ;
        RECT  0.695 0.380 0.865 0.555 ;
        RECT  0.470 0.750 0.660 0.960 ;
        RECT  0.400 0.750 0.470 1.180 ;
        RECT  0.350 0.840 0.400 1.180 ;
        RECT  0.255 1.060 0.350 1.180 ;
        RECT  0.135 1.060 0.255 1.555 ;
        RECT  0.085 1.385 0.135 1.555 ;
    END
END SDFFRQXLAD
MACRO SDFFRX1AD
    CLASS CORE ;
    FOREIGN SDFFRX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.865 1.665 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.705 0.430 1.935 ;
        END
        AntennaGateArea 0.108 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.545 0.990 6.665 1.250 ;
        RECT  6.160 0.990 6.545 1.110 ;
        RECT  6.040 0.440 6.160 1.110 ;
        RECT  5.450 0.440 6.040 0.560 ;
        RECT  5.330 0.440 5.450 0.655 ;
        RECT  4.810 0.535 5.330 0.655 ;
        RECT  4.690 0.380 4.810 0.655 ;
        RECT  3.170 0.380 4.690 0.500 ;
        RECT  3.050 0.380 3.170 0.540 ;
        RECT  2.450 0.420 3.050 0.540 ;
        RECT  2.330 0.420 2.450 0.980 ;
        RECT  2.170 0.860 2.330 0.980 ;
        RECT  2.030 0.860 2.170 1.375 ;
        RECT  2.025 1.255 2.030 1.375 ;
        RECT  1.855 1.255 2.025 1.535 ;
        END
        AntennaGateArea 0.123 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.350 0.680 7.530 1.600 ;
        END
        AntennaDiffArea 0.207 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.170 0.660 8.330 1.920 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.110 0.870 1.450 ;
        END
        AntennaGateArea 0.065 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.100 2.575 1.375 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.925 -0.210 8.400 0.210 ;
        RECT  7.755 -0.210 7.925 0.895 ;
        RECT  6.555 -0.210 7.755 0.210 ;
        RECT  6.295 -0.210 6.555 0.815 ;
        RECT  5.210 -0.210 6.295 0.210 ;
        RECT  4.950 -0.210 5.210 0.415 ;
        RECT  2.940 -0.210 4.950 0.210 ;
        RECT  2.420 -0.210 2.940 0.300 ;
        RECT  0.230 -0.210 2.420 0.210 ;
        RECT  0.110 -0.210 0.230 0.940 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.935 2.310 8.400 2.730 ;
        RECT  7.765 1.985 7.935 2.730 ;
        RECT  7.205 2.310 7.765 2.730 ;
        RECT  7.035 2.020 7.205 2.730 ;
        RECT  6.535 2.310 7.035 2.730 ;
        RECT  6.365 2.020 6.535 2.730 ;
        RECT  4.525 2.310 6.365 2.730 ;
        RECT  4.265 2.095 4.525 2.730 ;
        RECT  2.860 2.310 4.265 2.730 ;
        RECT  2.600 2.220 2.860 2.730 ;
        RECT  1.765 2.310 2.600 2.730 ;
        RECT  1.595 2.175 1.765 2.730 ;
        RECT  0.600 2.310 1.595 2.730 ;
        RECT  0.340 2.055 0.600 2.730 ;
        RECT  0.000 2.310 0.340 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.400 2.520 ;
        LAYER M1 ;
        RECT  7.930 1.020 8.050 1.865 ;
        RECT  7.215 1.745 7.930 1.865 ;
        RECT  7.095 0.625 7.215 1.865 ;
        RECT  7.005 0.625 7.095 0.885 ;
        RECT  6.240 1.615 7.095 1.735 ;
        RECT  6.855 1.125 6.975 1.490 ;
        RECT  5.780 1.370 6.855 1.490 ;
        RECT  6.120 1.615 6.240 2.115 ;
        RECT  5.830 2.070 5.970 2.190 ;
        RECT  5.780 0.695 5.920 0.815 ;
        RECT  5.710 1.925 5.830 2.190 ;
        RECT  5.660 0.695 5.780 1.805 ;
        RECT  5.060 1.925 5.710 2.045 ;
        RECT  5.620 1.545 5.660 1.805 ;
        RECT  5.310 0.790 5.455 1.805 ;
        RECT  5.300 1.270 5.310 1.805 ;
        RECT  4.640 1.270 5.300 1.390 ;
        RECT  5.260 1.545 5.300 1.805 ;
        RECT  4.940 1.585 5.060 2.045 ;
        RECT  4.400 1.585 4.940 1.705 ;
        RECT  4.700 1.855 4.820 2.120 ;
        RECT  4.160 1.855 4.700 1.975 ;
        RECT  4.520 1.205 4.640 1.465 ;
        RECT  4.280 0.620 4.400 1.705 ;
        RECT  3.540 0.620 4.280 0.740 ;
        RECT  4.040 0.890 4.160 1.975 ;
        RECT  3.760 1.855 4.040 1.975 ;
        RECT  3.715 0.890 3.835 1.735 ;
        RECT  3.580 1.855 3.760 2.100 ;
        RECT  3.660 0.890 3.715 1.150 ;
        RECT  3.460 1.615 3.715 1.735 ;
        RECT  1.930 1.980 3.580 2.100 ;
        RECT  3.540 1.235 3.575 1.495 ;
        RECT  3.420 0.620 3.540 1.495 ;
        RECT  3.245 1.615 3.460 1.860 ;
        RECT  3.340 0.620 3.420 0.740 ;
        RECT  3.105 1.315 3.420 1.495 ;
        RECT  3.180 0.885 3.300 1.145 ;
        RECT  1.350 1.740 3.245 1.860 ;
        RECT  2.815 1.025 3.180 1.145 ;
        RECT  2.935 1.315 3.105 1.560 ;
        RECT  2.815 0.660 2.880 0.780 ;
        RECT  2.695 0.660 2.815 1.615 ;
        RECT  2.620 0.660 2.695 0.780 ;
        RECT  2.220 1.495 2.695 1.615 ;
        RECT  1.955 0.380 2.125 0.695 ;
        RECT  0.650 0.380 1.955 0.500 ;
        RECT  1.350 0.620 1.540 0.740 ;
        RECT  1.230 0.620 1.350 1.860 ;
        RECT  1.025 1.660 1.230 1.860 ;
        RECT  0.990 0.840 1.110 1.360 ;
        RECT  0.660 0.840 0.990 0.960 ;
        RECT  0.470 0.750 0.660 0.960 ;
        RECT  0.400 0.750 0.470 1.180 ;
        RECT  0.350 0.840 0.400 1.180 ;
        RECT  0.255 1.060 0.350 1.180 ;
        RECT  0.135 1.060 0.255 1.555 ;
        RECT  0.085 1.385 0.135 1.555 ;
    END
END SDFFRX1AD
MACRO SDFFRX2AD
    CLASS CORE ;
    FOREIGN SDFFRX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.660 0.865 1.890 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.705 0.355 2.020 ;
        RECT  0.070 1.705 0.185 1.935 ;
        END
        AntennaGateArea 0.105 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.435 0.335 6.605 0.535 ;
        RECT  5.250 0.380 6.435 0.500 ;
        RECT  5.130 0.380 5.250 0.785 ;
        RECT  5.080 0.665 5.130 0.785 ;
        RECT  4.820 0.665 5.080 1.115 ;
        RECT  4.725 0.665 4.820 0.785 ;
        RECT  4.605 0.380 4.725 0.785 ;
        RECT  3.155 0.380 4.605 0.500 ;
        RECT  3.035 0.380 3.155 0.540 ;
        RECT  2.450 0.420 3.035 0.540 ;
        RECT  2.330 0.420 2.450 1.025 ;
        RECT  2.140 0.905 2.330 1.025 ;
        RECT  2.020 0.905 2.140 1.620 ;
        END
        AntennaGateArea 0.13 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.520 0.385 7.585 0.815 ;
        RECT  7.520 1.375 7.585 1.545 ;
        RECT  7.350 0.385 7.520 1.545 ;
        END
        AntennaDiffArea 0.373 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.190 0.340 8.330 2.030 ;
        RECT  8.160 0.340 8.190 0.860 ;
        RECT  8.160 1.510 8.190 2.030 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.605 1.110 0.910 1.375 ;
        END
        AntennaGateArea 0.064 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.580 1.020 2.700 1.375 ;
        RECT  2.310 1.145 2.580 1.375 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.945 -0.210 8.400 0.210 ;
        RECT  7.775 -0.210 7.945 0.815 ;
        RECT  6.845 -0.210 7.775 0.210 ;
        RECT  6.725 -0.210 6.845 0.810 ;
        RECT  5.010 -0.210 6.725 0.210 ;
        RECT  6.270 0.690 6.725 0.810 ;
        RECT  4.890 -0.210 5.010 0.460 ;
        RECT  2.925 -0.210 4.890 0.210 ;
        RECT  2.405 -0.210 2.925 0.300 ;
        RECT  0.230 -0.210 2.405 0.210 ;
        RECT  0.110 -0.210 0.230 0.940 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.945 2.310 8.400 2.730 ;
        RECT  7.775 1.945 7.945 2.730 ;
        RECT  7.245 2.310 7.775 2.730 ;
        RECT  7.075 1.920 7.245 2.730 ;
        RECT  6.530 2.310 7.075 2.730 ;
        RECT  6.270 1.595 6.530 2.730 ;
        RECT  5.010 2.310 6.270 2.730 ;
        RECT  4.840 1.780 5.010 2.730 ;
        RECT  4.480 2.310 4.840 2.730 ;
        RECT  4.220 2.130 4.480 2.730 ;
        RECT  2.900 2.310 4.220 2.730 ;
        RECT  2.640 2.220 2.900 2.730 ;
        RECT  1.960 2.310 2.640 2.730 ;
        RECT  1.700 1.980 1.960 2.730 ;
        RECT  0.645 2.310 1.700 2.730 ;
        RECT  0.475 1.505 0.645 2.730 ;
        RECT  0.000 2.310 0.475 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.400 2.520 ;
        LAYER M1 ;
        RECT  7.890 1.020 8.010 1.785 ;
        RECT  7.215 1.665 7.890 1.785 ;
        RECT  7.095 0.935 7.215 1.785 ;
        RECT  7.085 0.935 7.095 1.055 ;
        RECT  6.910 1.665 7.095 1.785 ;
        RECT  6.965 0.620 7.085 1.055 ;
        RECT  6.805 1.175 6.975 1.420 ;
        RECT  6.410 0.935 6.965 1.055 ;
        RECT  6.650 1.595 6.910 1.785 ;
        RECT  5.875 1.300 6.805 1.420 ;
        RECT  6.150 0.935 6.410 1.140 ;
        RECT  5.875 1.965 6.135 2.190 ;
        RECT  5.755 0.665 5.875 1.740 ;
        RECT  5.250 1.965 5.875 2.085 ;
        RECT  5.705 0.665 5.755 0.835 ;
        RECT  5.705 1.570 5.755 1.740 ;
        RECT  5.370 0.620 5.490 1.845 ;
        RECT  4.605 1.295 5.370 1.415 ;
        RECT  5.130 1.540 5.250 2.085 ;
        RECT  4.485 1.540 5.130 1.660 ;
        RECT  4.600 1.810 4.720 2.190 ;
        RECT  4.240 1.810 4.600 1.930 ;
        RECT  4.365 0.620 4.485 1.660 ;
        RECT  3.600 0.620 4.365 0.740 ;
        RECT  4.120 0.860 4.240 1.930 ;
        RECT  3.910 1.810 4.120 1.930 ;
        RECT  3.860 1.730 3.910 1.930 ;
        RECT  3.840 0.860 3.880 1.120 ;
        RECT  3.740 1.730 3.860 2.100 ;
        RECT  3.720 0.860 3.840 1.610 ;
        RECT  2.080 1.980 3.740 2.100 ;
        RECT  3.595 1.490 3.720 1.610 ;
        RECT  3.480 0.620 3.600 1.370 ;
        RECT  3.475 1.490 3.595 1.860 ;
        RECT  3.270 0.660 3.480 0.780 ;
        RECT  3.220 1.250 3.480 1.370 ;
        RECT  1.530 1.740 3.475 1.860 ;
        RECT  2.955 0.945 3.295 1.115 ;
        RECT  3.100 1.250 3.220 1.605 ;
        RECT  2.835 0.660 2.955 1.615 ;
        RECT  2.600 0.660 2.835 0.780 ;
        RECT  2.360 1.495 2.835 1.615 ;
        RECT  2.100 0.600 2.150 0.770 ;
        RECT  1.980 0.380 2.100 0.770 ;
        RECT  0.895 0.380 1.980 0.500 ;
        RECT  1.530 0.625 1.580 0.745 ;
        RECT  1.410 0.625 1.530 1.860 ;
        RECT  1.320 0.625 1.410 0.745 ;
        RECT  1.105 1.665 1.410 1.860 ;
        RECT  1.150 1.155 1.290 1.275 ;
        RECT  1.030 0.840 1.150 1.275 ;
        RECT  0.615 0.840 1.030 0.960 ;
        RECT  0.725 0.380 0.895 0.555 ;
        RECT  0.480 0.725 0.615 0.960 ;
        RECT  0.445 0.725 0.480 1.180 ;
        RECT  0.360 0.840 0.445 1.180 ;
        RECT  0.255 1.060 0.360 1.180 ;
        RECT  0.135 1.060 0.255 1.555 ;
        RECT  0.085 1.385 0.135 1.555 ;
    END
END SDFFRX2AD
MACRO SDFFRX4AD
    CLASS CORE ;
    FOREIGN SDFFRX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.865 1.945 1.300 ;
        END
        AntennaGateArea 0.06 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.185 1.705 0.355 2.020 ;
        RECT  0.070 1.705 0.185 1.935 ;
        END
        AntennaGateArea 0.142 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.170 0.775 6.700 0.895 ;
        RECT  6.050 0.380 6.170 0.895 ;
        RECT  5.280 0.380 6.050 0.500 ;
        RECT  5.160 0.380 5.280 0.705 ;
        RECT  5.090 0.585 5.160 0.705 ;
        RECT  5.040 0.585 5.090 1.020 ;
        RECT  4.920 0.585 5.040 1.200 ;
        RECT  4.830 0.585 4.920 1.020 ;
        RECT  4.800 0.585 4.830 0.705 ;
        RECT  4.680 0.380 4.800 0.705 ;
        RECT  3.155 0.380 4.680 0.500 ;
        RECT  3.035 0.380 3.155 0.540 ;
        RECT  2.465 0.420 3.035 0.540 ;
        RECT  2.345 0.420 2.465 1.265 ;
        RECT  2.220 1.145 2.345 1.265 ;
        RECT  2.100 1.145 2.220 1.655 ;
        RECT  1.960 1.535 2.100 1.655 ;
        END
        AntennaGateArea 0.191 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.625 0.385 7.795 1.545 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.540 0.975 8.610 1.515 ;
        RECT  8.370 0.340 8.540 2.030 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.605 1.020 0.910 1.375 ;
        END
        AntennaGateArea 0.108 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.920 2.750 1.375 ;
        END
        AntennaGateArea 0.114 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.875 -0.210 8.960 0.210 ;
        RECT  8.705 -0.210 8.875 0.815 ;
        RECT  8.155 -0.210 8.705 0.210 ;
        RECT  7.985 -0.210 8.155 0.815 ;
        RECT  7.410 -0.210 7.985 0.210 ;
        RECT  7.290 -0.210 7.410 0.930 ;
        RECT  6.515 -0.210 7.290 0.210 ;
        RECT  6.515 0.495 6.580 0.615 ;
        RECT  6.395 -0.210 6.515 0.615 ;
        RECT  5.040 -0.210 6.395 0.210 ;
        RECT  6.320 0.495 6.395 0.615 ;
        RECT  4.920 -0.210 5.040 0.460 ;
        RECT  3.240 -0.210 4.920 0.210 ;
        RECT  2.980 -0.210 3.240 0.250 ;
        RECT  2.655 -0.210 2.980 0.210 ;
        RECT  2.395 -0.210 2.655 0.250 ;
        RECT  0.230 -0.210 2.395 0.210 ;
        RECT  0.110 -0.210 0.230 0.940 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.875 2.310 8.960 2.730 ;
        RECT  8.705 1.670 8.875 2.730 ;
        RECT  8.155 2.310 8.705 2.730 ;
        RECT  7.985 1.945 8.155 2.730 ;
        RECT  7.395 2.310 7.985 2.730 ;
        RECT  7.225 1.920 7.395 2.730 ;
        RECT  6.535 2.310 7.225 2.730 ;
        RECT  6.365 1.575 6.535 2.730 ;
        RECT  5.060 2.310 6.365 2.730 ;
        RECT  4.890 1.820 5.060 2.730 ;
        RECT  2.990 2.310 4.890 2.730 ;
        RECT  2.730 2.260 2.990 2.730 ;
        RECT  1.960 2.310 2.730 2.730 ;
        RECT  1.700 2.020 1.960 2.730 ;
        RECT  0.645 2.310 1.700 2.730 ;
        RECT  0.475 1.505 0.645 2.730 ;
        RECT  0.000 2.310 0.475 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.960 2.520 ;
        LAYER M1 ;
        RECT  8.100 1.020 8.220 1.785 ;
        RECT  7.420 1.665 8.100 1.785 ;
        RECT  7.300 1.075 7.420 1.785 ;
        RECT  7.140 1.075 7.300 1.195 ;
        RECT  6.965 1.665 7.300 1.785 ;
        RECT  7.020 0.330 7.140 1.195 ;
        RECT  5.930 1.315 7.085 1.435 ;
        RECT  6.200 1.075 7.020 1.195 ;
        RECT  6.705 1.600 6.965 1.785 ;
        RECT  5.920 1.965 6.190 2.190 ;
        RECT  5.925 1.315 5.930 1.730 ;
        RECT  5.905 1.315 5.925 1.745 ;
        RECT  5.300 1.965 5.920 2.085 ;
        RECT  5.785 0.665 5.905 1.745 ;
        RECT  5.735 0.665 5.785 0.835 ;
        RECT  5.755 1.575 5.785 1.745 ;
        RECT  5.420 0.620 5.540 1.845 ;
        RECT  5.400 0.620 5.420 1.460 ;
        RECT  4.630 1.340 5.400 1.460 ;
        RECT  5.180 1.580 5.300 2.085 ;
        RECT  4.490 1.580 5.180 1.700 ;
        RECT  4.645 1.825 4.765 2.190 ;
        RECT  4.250 1.825 4.645 1.945 ;
        RECT  4.370 0.620 4.490 1.700 ;
        RECT  3.600 0.620 4.370 0.740 ;
        RECT  4.130 0.860 4.250 1.945 ;
        RECT  3.985 1.730 4.130 1.945 ;
        RECT  3.865 1.730 3.985 2.140 ;
        RECT  3.760 0.860 3.880 1.610 ;
        RECT  2.080 2.020 3.865 2.140 ;
        RECT  3.720 1.490 3.760 1.610 ;
        RECT  3.600 1.490 3.720 1.900 ;
        RECT  3.480 0.620 3.600 1.370 ;
        RECT  1.630 1.780 3.600 1.900 ;
        RECT  3.335 0.620 3.480 0.805 ;
        RECT  3.370 1.250 3.480 1.370 ;
        RECT  3.250 1.250 3.370 1.660 ;
        RECT  2.990 0.945 3.295 1.115 ;
        RECT  3.110 1.540 3.250 1.660 ;
        RECT  2.870 0.660 2.990 1.615 ;
        RECT  2.600 0.660 2.870 0.780 ;
        RECT  2.350 1.495 2.870 1.615 ;
        RECT  2.010 0.380 2.180 0.720 ;
        RECT  0.955 0.380 2.010 0.500 ;
        RECT  1.510 0.620 1.630 1.900 ;
        RECT  1.350 0.620 1.510 0.740 ;
        RECT  1.105 1.515 1.510 1.710 ;
        RECT  1.270 0.995 1.390 1.255 ;
        RECT  1.230 0.995 1.270 1.115 ;
        RECT  1.110 0.775 1.230 1.115 ;
        RECT  0.615 0.775 1.110 0.895 ;
        RECT  0.785 0.380 0.955 0.655 ;
        RECT  0.470 0.725 0.615 0.895 ;
        RECT  0.445 0.725 0.470 1.180 ;
        RECT  0.350 0.775 0.445 1.180 ;
        RECT  0.255 1.060 0.350 1.180 ;
        RECT  0.135 1.060 0.255 1.555 ;
        RECT  0.085 1.385 0.135 1.555 ;
    END
END SDFFRX4AD
MACRO SDFFRXLAD
    CLASS CORE ;
    FOREIGN SDFFRXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.865 1.665 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.705 0.430 1.935 ;
        END
        AntennaGateArea 0.106 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.545 0.990 6.665 1.250 ;
        RECT  6.160 0.990 6.545 1.110 ;
        RECT  6.040 0.440 6.160 1.110 ;
        RECT  5.450 0.440 6.040 0.560 ;
        RECT  5.330 0.440 5.450 0.655 ;
        RECT  4.810 0.535 5.330 0.655 ;
        RECT  4.690 0.380 4.810 0.655 ;
        RECT  3.170 0.380 4.690 0.500 ;
        RECT  3.050 0.380 3.170 0.540 ;
        RECT  2.450 0.420 3.050 0.540 ;
        RECT  2.330 0.420 2.450 0.980 ;
        RECT  2.170 0.860 2.330 0.980 ;
        RECT  2.030 0.860 2.170 1.375 ;
        RECT  2.025 1.255 2.030 1.375 ;
        RECT  1.855 1.255 2.025 1.535 ;
        END
        AntennaGateArea 0.124 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.350 0.680 7.530 1.600 ;
        END
        AntennaDiffArea 0.14 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.170 0.690 8.330 1.695 ;
        END
        AntennaDiffArea 0.138 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.110 0.870 1.450 ;
        END
        AntennaGateArea 0.065 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.100 2.575 1.375 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.970 -0.210 8.400 0.210 ;
        RECT  7.710 -0.210 7.970 0.880 ;
        RECT  6.555 -0.210 7.710 0.210 ;
        RECT  6.295 -0.210 6.555 0.815 ;
        RECT  5.210 -0.210 6.295 0.210 ;
        RECT  4.950 -0.210 5.210 0.415 ;
        RECT  2.940 -0.210 4.950 0.210 ;
        RECT  2.420 -0.210 2.940 0.300 ;
        RECT  0.230 -0.210 2.420 0.210 ;
        RECT  0.110 -0.210 0.230 0.940 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.935 2.310 8.400 2.730 ;
        RECT  7.765 1.985 7.935 2.730 ;
        RECT  7.205 2.310 7.765 2.730 ;
        RECT  7.035 2.020 7.205 2.730 ;
        RECT  6.535 2.310 7.035 2.730 ;
        RECT  6.365 2.020 6.535 2.730 ;
        RECT  4.525 2.310 6.365 2.730 ;
        RECT  4.265 2.095 4.525 2.730 ;
        RECT  2.860 2.310 4.265 2.730 ;
        RECT  2.600 2.220 2.860 2.730 ;
        RECT  1.765 2.310 2.600 2.730 ;
        RECT  1.595 2.175 1.765 2.730 ;
        RECT  0.600 2.310 1.595 2.730 ;
        RECT  0.340 2.055 0.600 2.730 ;
        RECT  0.000 2.310 0.340 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.400 2.520 ;
        LAYER M1 ;
        RECT  7.930 1.020 8.050 1.865 ;
        RECT  7.215 1.745 7.930 1.865 ;
        RECT  7.095 0.625 7.215 1.865 ;
        RECT  7.005 0.625 7.095 0.885 ;
        RECT  6.240 1.615 7.095 1.735 ;
        RECT  6.855 1.125 6.975 1.490 ;
        RECT  5.780 1.370 6.855 1.490 ;
        RECT  6.120 1.615 6.240 2.115 ;
        RECT  5.830 2.070 5.970 2.190 ;
        RECT  5.780 0.695 5.920 0.815 ;
        RECT  5.710 1.925 5.830 2.190 ;
        RECT  5.660 0.695 5.780 1.805 ;
        RECT  5.060 1.925 5.710 2.045 ;
        RECT  5.620 1.545 5.660 1.805 ;
        RECT  5.310 0.790 5.455 1.805 ;
        RECT  5.300 1.270 5.310 1.805 ;
        RECT  4.640 1.270 5.300 1.390 ;
        RECT  5.260 1.545 5.300 1.805 ;
        RECT  4.940 1.585 5.060 2.045 ;
        RECT  4.400 1.585 4.940 1.705 ;
        RECT  4.700 1.855 4.820 2.120 ;
        RECT  4.160 1.855 4.700 1.975 ;
        RECT  4.520 1.205 4.640 1.465 ;
        RECT  4.280 0.620 4.400 1.705 ;
        RECT  3.540 0.620 4.280 0.740 ;
        RECT  4.040 0.890 4.160 1.975 ;
        RECT  3.760 1.855 4.040 1.975 ;
        RECT  3.715 0.890 3.835 1.735 ;
        RECT  3.580 1.855 3.760 2.100 ;
        RECT  3.660 0.890 3.715 1.150 ;
        RECT  3.460 1.615 3.715 1.735 ;
        RECT  1.930 1.980 3.580 2.100 ;
        RECT  3.540 1.235 3.575 1.495 ;
        RECT  3.420 0.620 3.540 1.495 ;
        RECT  3.245 1.615 3.460 1.860 ;
        RECT  3.340 0.620 3.420 0.740 ;
        RECT  3.105 1.315 3.420 1.495 ;
        RECT  3.180 0.885 3.300 1.145 ;
        RECT  1.350 1.740 3.245 1.860 ;
        RECT  2.815 1.025 3.180 1.145 ;
        RECT  2.935 1.315 3.105 1.560 ;
        RECT  2.815 0.660 2.880 0.780 ;
        RECT  2.695 0.660 2.815 1.615 ;
        RECT  2.620 0.660 2.695 0.780 ;
        RECT  2.220 1.495 2.695 1.615 ;
        RECT  1.955 0.380 2.125 0.695 ;
        RECT  0.650 0.380 1.955 0.500 ;
        RECT  1.350 0.620 1.540 0.740 ;
        RECT  1.230 0.620 1.350 1.860 ;
        RECT  1.025 1.660 1.230 1.860 ;
        RECT  0.990 0.840 1.110 1.360 ;
        RECT  0.660 0.840 0.990 0.960 ;
        RECT  0.470 0.750 0.660 0.960 ;
        RECT  0.400 0.750 0.470 1.180 ;
        RECT  0.350 0.840 0.400 1.180 ;
        RECT  0.255 1.060 0.350 1.180 ;
        RECT  0.135 1.060 0.255 1.555 ;
        RECT  0.085 1.385 0.135 1.555 ;
    END
END SDFFRXLAD
MACRO SDFFSHQX1AD
    CLASS CORE ;
    FOREIGN SDFFSHQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.675 1.190 4.735 1.330 ;
        RECT  4.350 0.960 4.675 1.330 ;
        RECT  4.285 0.960 4.350 1.220 ;
        END
        AntennaGateArea 0.109 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.625 0.800 3.850 1.095 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.905 1.325 3.025 1.660 ;
        RECT  2.370 1.540 2.905 1.660 ;
        RECT  2.250 1.245 2.370 1.660 ;
        RECT  2.215 1.245 2.250 1.365 ;
        RECT  2.120 1.190 2.215 1.365 ;
        RECT  1.985 1.035 2.120 1.365 ;
        END
        AntennaGateArea 0.101 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.290 0.600 9.450 1.930 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.320 0.865 2.495 1.125 ;
        RECT  2.240 0.865 2.320 1.050 ;
        END
        AntennaGateArea 0.056 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.000 0.530 1.375 ;
        END
        AntennaGateArea 0.114 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.055 -0.210 9.520 0.210 ;
        RECT  8.885 -0.210 9.055 0.335 ;
        RECT  8.225 -0.210 8.885 0.210 ;
        RECT  7.965 -0.210 8.225 0.330 ;
        RECT  6.380 -0.210 7.965 0.210 ;
        RECT  6.210 -0.210 6.380 0.260 ;
        RECT  4.330 -0.210 6.210 0.210 ;
        RECT  3.810 -0.210 4.330 0.260 ;
        RECT  2.265 -0.210 3.810 0.210 ;
        RECT  2.095 -0.210 2.265 0.260 ;
        RECT  1.165 -0.210 2.095 0.210 ;
        RECT  0.995 -0.210 1.165 0.375 ;
        RECT  0.635 -0.210 0.995 0.210 ;
        RECT  0.465 -0.210 0.635 0.375 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.010 2.310 9.520 2.730 ;
        RECT  8.570 1.965 9.010 2.730 ;
        RECT  6.850 2.310 8.570 2.730 ;
        RECT  6.680 1.925 6.850 2.730 ;
        RECT  5.715 2.310 6.680 2.730 ;
        RECT  5.595 2.150 5.715 2.730 ;
        RECT  4.455 2.310 5.595 2.730 ;
        RECT  4.285 2.145 4.455 2.730 ;
        RECT  2.385 2.310 4.285 2.730 ;
        RECT  2.215 2.260 2.385 2.730 ;
        RECT  1.835 2.310 2.215 2.730 ;
        RECT  1.665 2.260 1.835 2.730 ;
        RECT  0.555 2.310 1.665 2.730 ;
        RECT  0.385 1.915 0.555 2.730 ;
        RECT  0.000 2.310 0.385 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.520 2.520 ;
        LAYER M1 ;
        RECT  8.925 0.455 9.045 1.840 ;
        RECT  8.560 0.455 8.925 0.575 ;
        RECT  8.395 1.720 8.925 1.840 ;
        RECT  8.535 0.695 8.705 1.545 ;
        RECT  8.390 0.355 8.560 0.575 ;
        RECT  8.275 1.070 8.535 1.240 ;
        RECT  8.275 1.720 8.395 2.045 ;
        RECT  7.405 0.455 8.390 0.575 ;
        RECT  8.155 0.755 8.365 0.875 ;
        RECT  7.445 1.925 8.275 2.045 ;
        RECT  8.035 0.755 8.155 1.805 ;
        RECT  6.435 1.685 8.035 1.805 ;
        RECT  7.735 0.925 7.855 1.565 ;
        RECT  7.165 0.925 7.735 1.045 ;
        RECT  7.285 0.420 7.405 0.680 ;
        RECT  6.885 1.405 7.325 1.565 ;
        RECT  7.045 0.380 7.165 1.045 ;
        RECT  5.795 0.380 7.045 0.500 ;
        RECT  6.765 0.670 6.885 1.565 ;
        RECT  6.555 1.375 6.765 1.565 ;
        RECT  6.525 0.620 6.645 1.255 ;
        RECT  4.165 0.620 6.525 0.740 ;
        RECT  6.435 1.135 6.525 1.255 ;
        RECT  6.315 1.135 6.435 1.805 ;
        RECT  5.645 0.895 6.405 1.015 ;
        RECT  6.125 2.020 6.385 2.190 ;
        RECT  6.075 1.490 6.195 1.900 ;
        RECT  5.955 2.020 6.125 2.140 ;
        RECT  5.505 1.490 6.075 1.610 ;
        RECT  5.835 1.880 5.955 2.140 ;
        RECT  5.055 1.880 5.835 2.000 ;
        RECT  5.535 0.335 5.795 0.500 ;
        RECT  5.505 0.860 5.645 1.015 ;
        RECT  1.550 0.380 5.535 0.500 ;
        RECT  5.385 0.860 5.505 1.610 ;
        RECT  5.305 1.490 5.385 1.610 ;
        RECT  5.185 1.490 5.305 1.750 ;
        RECT  5.055 0.935 5.100 1.055 ;
        RECT  4.935 0.935 5.055 2.025 ;
        RECT  4.840 0.935 4.935 1.055 ;
        RECT  4.165 1.905 4.935 2.025 ;
        RECT  4.610 1.615 4.780 1.785 ;
        RECT  3.925 1.665 4.610 1.785 ;
        RECT  4.165 1.375 4.230 1.545 ;
        RECT  4.045 0.620 4.165 1.545 ;
        RECT  4.045 1.905 4.165 2.140 ;
        RECT  3.970 0.620 4.045 0.740 ;
        RECT  1.890 2.020 4.045 2.140 ;
        RECT  3.805 1.215 3.925 1.900 ;
        RECT  3.505 1.215 3.805 1.335 ;
        RECT  3.385 1.780 3.805 1.900 ;
        RECT  3.265 1.475 3.685 1.645 ;
        RECT  3.385 0.625 3.505 1.335 ;
        RECT  2.880 0.625 3.385 0.745 ;
        RECT  3.145 1.005 3.265 1.900 ;
        RECT  3.000 1.005 3.145 1.125 ;
        RECT  2.130 1.780 3.145 1.900 ;
        RECT  2.880 0.865 3.000 1.125 ;
        RECT  2.735 1.250 2.785 1.420 ;
        RECT  2.615 0.625 2.735 1.420 ;
        RECT  2.430 0.625 2.615 0.745 ;
        RECT  2.010 1.485 2.130 1.900 ;
        RECT  1.790 1.485 2.010 1.605 ;
        RECT  1.790 0.625 1.980 0.745 ;
        RECT  1.770 1.875 1.890 2.140 ;
        RECT  1.670 0.625 1.790 1.605 ;
        RECT  1.160 1.875 1.770 1.995 ;
        RECT  1.430 0.335 1.550 1.520 ;
        RECT  1.010 1.400 1.430 1.520 ;
        RECT  1.190 0.495 1.310 1.195 ;
        RECT  0.230 0.495 1.190 0.615 ;
        RECT  1.040 1.670 1.160 1.995 ;
        RECT  0.770 1.670 1.040 1.790 ;
        RECT  0.890 1.020 1.010 1.520 ;
        RECT  0.770 0.760 0.980 0.880 ;
        RECT  0.650 0.760 0.770 1.790 ;
        RECT  0.110 0.495 0.230 1.590 ;
    END
END SDFFSHQX1AD
MACRO SDFFSHQX2AD
    CLASS CORE ;
    FOREIGN SDFFSHQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.350 0.980 4.740 1.330 ;
        RECT  4.285 0.980 4.350 1.240 ;
        END
        AntennaGateArea 0.135 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.625 0.800 3.850 1.095 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.905 1.325 3.025 1.660 ;
        RECT  2.370 1.540 2.905 1.660 ;
        RECT  2.250 1.245 2.370 1.660 ;
        RECT  2.215 1.245 2.250 1.365 ;
        RECT  2.120 1.190 2.215 1.365 ;
        RECT  1.985 1.035 2.120 1.365 ;
        END
        AntennaGateArea 0.118 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.290 0.600 9.450 2.190 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.320 0.865 2.495 1.125 ;
        RECT  2.240 0.865 2.320 1.050 ;
        END
        AntennaGateArea 0.086 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.000 0.530 1.375 ;
        END
        AntennaGateArea 0.121 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.005 -0.210 9.520 0.210 ;
        RECT  8.835 -0.210 9.005 0.335 ;
        RECT  8.225 -0.210 8.835 0.210 ;
        RECT  7.965 -0.210 8.225 0.330 ;
        RECT  6.450 -0.210 7.965 0.210 ;
        RECT  6.020 -0.210 6.450 0.260 ;
        RECT  4.330 -0.210 6.020 0.210 ;
        RECT  3.810 -0.210 4.330 0.260 ;
        RECT  2.265 -0.210 3.810 0.210 ;
        RECT  2.095 -0.210 2.265 0.260 ;
        RECT  1.165 -0.210 2.095 0.210 ;
        RECT  0.995 -0.210 1.165 0.375 ;
        RECT  0.635 -0.210 0.995 0.210 ;
        RECT  0.465 -0.210 0.635 0.375 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.005 2.310 9.520 2.730 ;
        RECT  8.575 1.965 9.005 2.730 ;
        RECT  6.850 2.310 8.575 2.730 ;
        RECT  6.680 1.925 6.850 2.730 ;
        RECT  6.005 2.310 6.680 2.730 ;
        RECT  5.745 2.290 6.005 2.730 ;
        RECT  4.455 2.310 5.745 2.730 ;
        RECT  4.285 2.260 4.455 2.730 ;
        RECT  2.385 2.310 4.285 2.730 ;
        RECT  2.215 2.260 2.385 2.730 ;
        RECT  1.835 2.310 2.215 2.730 ;
        RECT  1.665 2.260 1.835 2.730 ;
        RECT  0.555 2.310 1.665 2.730 ;
        RECT  0.385 1.865 0.555 2.730 ;
        RECT  0.000 2.310 0.385 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.520 2.520 ;
        LAYER M1 ;
        RECT  8.925 0.455 9.045 1.840 ;
        RECT  8.560 0.455 8.925 0.575 ;
        RECT  8.395 1.720 8.925 1.840 ;
        RECT  8.535 0.695 8.705 1.545 ;
        RECT  8.390 0.355 8.560 0.575 ;
        RECT  8.275 1.070 8.535 1.240 ;
        RECT  8.275 1.720 8.395 2.045 ;
        RECT  7.405 0.455 8.390 0.575 ;
        RECT  8.155 0.755 8.365 0.875 ;
        RECT  7.445 1.925 8.275 2.045 ;
        RECT  8.035 0.755 8.155 1.805 ;
        RECT  6.435 1.685 8.035 1.805 ;
        RECT  7.735 0.925 7.855 1.565 ;
        RECT  7.165 0.925 7.735 1.045 ;
        RECT  7.285 0.455 7.405 0.715 ;
        RECT  6.905 1.405 7.325 1.565 ;
        RECT  7.045 0.380 7.165 1.045 ;
        RECT  5.795 0.380 7.045 0.500 ;
        RECT  6.735 0.620 6.905 1.565 ;
        RECT  6.555 1.375 6.735 1.565 ;
        RECT  6.495 0.620 6.615 1.255 ;
        RECT  4.165 0.620 6.495 0.740 ;
        RECT  6.435 1.135 6.495 1.255 ;
        RECT  6.315 1.135 6.435 1.805 ;
        RECT  6.125 2.020 6.385 2.190 ;
        RECT  5.645 0.895 6.375 1.015 ;
        RECT  6.075 1.490 6.195 1.900 ;
        RECT  5.955 2.020 6.125 2.140 ;
        RECT  5.505 1.490 6.075 1.610 ;
        RECT  5.835 1.880 5.955 2.140 ;
        RECT  5.055 1.880 5.835 2.000 ;
        RECT  5.535 0.335 5.795 0.500 ;
        RECT  5.505 0.860 5.645 1.015 ;
        RECT  1.550 0.380 5.535 0.500 ;
        RECT  5.385 0.860 5.505 1.610 ;
        RECT  5.330 1.490 5.385 1.610 ;
        RECT  5.160 1.490 5.330 1.745 ;
        RECT  5.030 1.880 5.055 2.140 ;
        RECT  4.910 0.960 5.030 2.140 ;
        RECT  1.890 2.020 4.910 2.140 ;
        RECT  4.610 1.730 4.780 1.900 ;
        RECT  3.925 1.780 4.610 1.900 ;
        RECT  4.165 1.375 4.230 1.545 ;
        RECT  4.045 0.620 4.165 1.545 ;
        RECT  3.970 0.620 4.045 0.740 ;
        RECT  3.805 1.215 3.925 1.900 ;
        RECT  3.505 1.215 3.805 1.335 ;
        RECT  3.385 1.780 3.805 1.900 ;
        RECT  3.265 1.475 3.685 1.645 ;
        RECT  3.385 0.625 3.505 1.335 ;
        RECT  2.880 0.625 3.385 0.745 ;
        RECT  3.145 1.005 3.265 1.900 ;
        RECT  3.000 1.005 3.145 1.125 ;
        RECT  2.130 1.780 3.145 1.900 ;
        RECT  2.880 0.865 3.000 1.125 ;
        RECT  2.735 1.250 2.785 1.420 ;
        RECT  2.615 0.625 2.735 1.420 ;
        RECT  2.430 0.625 2.615 0.745 ;
        RECT  2.010 1.485 2.130 1.900 ;
        RECT  1.790 1.485 2.010 1.605 ;
        RECT  1.790 0.625 1.980 0.745 ;
        RECT  1.770 1.875 1.890 2.140 ;
        RECT  1.670 0.625 1.790 1.605 ;
        RECT  1.160 1.875 1.770 1.995 ;
        RECT  1.430 0.335 1.550 1.520 ;
        RECT  1.010 1.400 1.430 1.520 ;
        RECT  1.190 0.495 1.310 1.195 ;
        RECT  0.230 0.495 1.190 0.615 ;
        RECT  1.040 1.670 1.160 1.995 ;
        RECT  0.770 1.670 1.040 1.790 ;
        RECT  0.890 1.020 1.010 1.520 ;
        RECT  0.770 0.755 0.980 0.875 ;
        RECT  0.650 0.755 0.770 1.790 ;
        RECT  0.110 0.495 0.230 1.600 ;
    END
END SDFFSHQX2AD
MACRO SDFFSHQX4AD
    CLASS CORE ;
    FOREIGN SDFFSHQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.495 0.960 4.885 1.375 ;
        END
        AntennaGateArea 0.156 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.520 1.150 3.895 1.330 ;
        END
        AntennaGateArea 0.055 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 1.245 3.130 1.660 ;
        RECT  1.890 1.540 3.010 1.660 ;
        RECT  1.750 1.105 1.890 1.660 ;
        RECT  1.585 1.105 1.750 1.535 ;
        END
        AntennaGateArea 0.146 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.035 1.005 11.130 1.515 ;
        RECT  10.865 0.415 11.035 2.120 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.865 2.625 1.150 ;
        END
        AntennaGateArea 0.135 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.325 1.025 0.530 1.445 ;
        END
        AntennaGateArea 0.192 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.395 -0.210 11.480 0.210 ;
        RECT  11.225 -0.210 11.395 0.845 ;
        RECT  10.675 -0.210 11.225 0.210 ;
        RECT  10.505 -0.210 10.675 0.845 ;
        RECT  9.445 -0.210 10.505 0.210 ;
        RECT  9.275 -0.210 9.445 0.325 ;
        RECT  7.740 -0.210 9.275 0.210 ;
        RECT  7.480 -0.210 7.740 0.630 ;
        RECT  6.840 -0.210 7.480 0.210 ;
        RECT  6.580 -0.210 6.840 0.500 ;
        RECT  5.020 -0.210 6.580 0.210 ;
        RECT  4.760 -0.210 5.020 0.230 ;
        RECT  4.520 -0.210 4.760 0.210 ;
        RECT  4.260 -0.210 4.520 0.230 ;
        RECT  3.920 -0.210 4.260 0.210 ;
        RECT  3.660 -0.210 3.920 0.255 ;
        RECT  2.290 -0.210 3.660 0.210 ;
        RECT  2.170 -0.210 2.290 0.500 ;
        RECT  1.490 -0.210 2.170 0.210 ;
        RECT  1.230 -0.210 1.490 0.230 ;
        RECT  0.680 -0.210 1.230 0.210 ;
        RECT  0.420 -0.210 0.680 0.230 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.395 2.310 11.480 2.730 ;
        RECT  11.225 1.635 11.395 2.730 ;
        RECT  10.570 2.310 11.225 2.730 ;
        RECT  10.140 1.960 10.570 2.730 ;
        RECT  8.090 2.310 10.140 2.730 ;
        RECT  7.920 1.910 8.090 2.730 ;
        RECT  7.280 2.310 7.920 2.730 ;
        RECT  7.110 1.910 7.280 2.730 ;
        RECT  6.315 2.310 7.110 2.730 ;
        RECT  6.055 2.190 6.315 2.730 ;
        RECT  4.785 2.310 6.055 2.730 ;
        RECT  4.615 2.260 4.785 2.730 ;
        RECT  4.335 2.310 4.615 2.730 ;
        RECT  4.165 2.260 4.335 2.730 ;
        RECT  2.625 2.310 4.165 2.730 ;
        RECT  2.365 2.290 2.625 2.730 ;
        RECT  1.595 2.310 2.365 2.730 ;
        RECT  1.335 2.260 1.595 2.730 ;
        RECT  0.600 2.310 1.335 2.730 ;
        RECT  0.430 2.075 0.600 2.730 ;
        RECT  0.000 2.310 0.430 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.480 2.520 ;
        LAYER M1 ;
        RECT  10.440 0.990 10.700 1.250 ;
        RECT  10.385 0.990 10.440 1.840 ;
        RECT  10.320 0.445 10.385 1.840 ;
        RECT  10.265 0.445 10.320 1.200 ;
        RECT  9.910 1.720 10.320 1.840 ;
        RECT  8.785 0.445 10.265 0.565 ;
        RECT  10.145 1.375 10.200 1.545 ;
        RECT  10.025 0.690 10.145 1.545 ;
        RECT  9.985 1.070 10.025 1.545 ;
        RECT  9.855 1.070 9.985 1.240 ;
        RECT  9.790 1.720 9.910 2.055 ;
        RECT  9.670 0.755 9.810 0.875 ;
        RECT  8.215 1.935 9.790 2.055 ;
        RECT  9.550 0.755 9.670 1.790 ;
        RECT  6.825 1.670 9.550 1.790 ;
        RECT  9.240 1.040 9.360 1.525 ;
        RECT  8.350 1.040 9.240 1.160 ;
        RECT  7.310 1.430 8.840 1.550 ;
        RECT  8.615 0.380 8.785 0.565 ;
        RECT  8.065 0.380 8.615 0.500 ;
        RECT  8.210 0.620 8.470 0.870 ;
        RECT  8.090 0.990 8.350 1.160 ;
        RECT  7.310 0.750 8.210 0.870 ;
        RECT  7.895 0.380 8.065 0.630 ;
        RECT  7.190 0.540 7.310 1.550 ;
        RECT  6.945 1.430 7.190 1.550 ;
        RECT  6.950 0.620 7.070 1.270 ;
        RECT  4.375 0.620 6.950 0.740 ;
        RECT  6.825 1.150 6.950 1.270 ;
        RECT  6.705 1.150 6.825 1.790 ;
        RECT  6.560 0.860 6.820 1.030 ;
        RECT  6.525 1.950 6.785 2.190 ;
        RECT  6.325 1.575 6.585 1.830 ;
        RECT  5.880 0.860 6.560 0.980 ;
        RECT  5.375 1.950 6.525 2.070 ;
        RECT  5.880 1.575 6.325 1.695 ;
        RECT  5.920 0.330 6.180 0.500 ;
        RECT  2.530 0.380 5.920 0.500 ;
        RECT  5.760 0.860 5.880 1.695 ;
        RECT  5.615 1.510 5.760 1.695 ;
        RECT  5.495 1.510 5.615 1.770 ;
        RECT  5.375 1.030 5.540 1.150 ;
        RECT  5.255 1.030 5.375 2.140 ;
        RECT  1.185 2.020 5.255 2.140 ;
        RECT  4.135 1.780 5.090 1.900 ;
        RECT  4.255 0.620 4.375 1.560 ;
        RECT  4.085 0.620 4.255 0.790 ;
        RECT  4.015 0.910 4.135 1.900 ;
        RECT  3.610 0.910 4.015 1.030 ;
        RECT  3.490 1.780 4.015 1.900 ;
        RECT  3.370 1.500 3.870 1.620 ;
        RECT  3.490 0.625 3.610 1.030 ;
        RECT  3.030 0.625 3.490 0.745 ;
        RECT  3.250 1.005 3.370 1.900 ;
        RECT  3.110 1.005 3.250 1.125 ;
        RECT  1.425 1.780 3.250 1.900 ;
        RECT  2.990 0.865 3.110 1.125 ;
        RECT  2.865 0.625 2.910 0.745 ;
        RECT  2.865 1.250 2.890 1.420 ;
        RECT  2.745 0.625 2.865 1.420 ;
        RECT  2.650 0.625 2.745 0.745 ;
        RECT  2.720 1.250 2.745 1.420 ;
        RECT  2.410 0.380 2.530 0.740 ;
        RECT  2.180 0.620 2.410 0.740 ;
        RECT  2.010 0.620 2.180 1.420 ;
        RECT  1.790 0.330 2.050 0.500 ;
        RECT  1.150 0.620 2.010 0.740 ;
        RECT  0.670 0.380 1.790 0.500 ;
        RECT  1.425 0.860 1.530 0.980 ;
        RECT  1.305 0.860 1.425 1.900 ;
        RECT  1.270 0.860 1.305 0.980 ;
        RECT  1.065 1.485 1.185 2.140 ;
        RECT  1.030 0.620 1.150 1.340 ;
        RECT  0.770 1.485 1.065 1.605 ;
        RECT  0.890 1.220 1.030 1.340 ;
        RECT  0.790 0.620 0.910 0.950 ;
        RECT  0.770 0.825 0.790 0.950 ;
        RECT  0.650 0.825 0.770 1.605 ;
        RECT  0.550 0.380 0.670 0.705 ;
        RECT  0.255 0.585 0.550 0.705 ;
        RECT  0.205 0.585 0.255 0.820 ;
        RECT  0.205 1.560 0.255 1.730 ;
        RECT  0.085 0.585 0.205 1.730 ;
    END
END SDFFSHQX4AD
MACRO SDFFSHQX8AD
    CLASS CORE ;
    FOREIGN SDFFSHQX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.495 0.960 4.885 1.375 ;
        END
        AntennaGateArea 0.166 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.520 1.150 3.895 1.330 ;
        END
        AntennaGateArea 0.103 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 1.245 3.130 1.660 ;
        RECT  1.890 1.540 3.010 1.660 ;
        RECT  1.750 1.105 1.890 1.660 ;
        RECT  1.585 1.105 1.750 1.535 ;
        END
        AntennaGateArea 0.167 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.585 0.370 11.755 2.170 ;
        RECT  11.035 1.005 11.585 1.515 ;
        RECT  10.850 0.370 11.035 2.170 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.865 2.625 1.150 ;
        END
        AntennaGateArea 0.135 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.325 0.995 0.530 1.375 ;
        END
        AntennaGateArea 0.256 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.115 -0.210 12.320 0.210 ;
        RECT  11.945 -0.210 12.115 0.800 ;
        RECT  11.395 -0.210 11.945 0.210 ;
        RECT  11.225 -0.210 11.395 0.800 ;
        RECT  10.675 -0.210 11.225 0.210 ;
        RECT  10.505 -0.210 10.675 0.800 ;
        RECT  9.445 -0.210 10.505 0.210 ;
        RECT  9.275 -0.210 9.445 0.325 ;
        RECT  7.740 -0.210 9.275 0.210 ;
        RECT  7.480 -0.210 7.740 0.630 ;
        RECT  6.840 -0.210 7.480 0.210 ;
        RECT  6.580 -0.210 6.840 0.500 ;
        RECT  5.020 -0.210 6.580 0.210 ;
        RECT  4.760 -0.210 5.020 0.240 ;
        RECT  4.520 -0.210 4.760 0.210 ;
        RECT  4.260 -0.210 4.520 0.240 ;
        RECT  3.920 -0.210 4.260 0.210 ;
        RECT  3.660 -0.210 3.920 0.255 ;
        RECT  2.290 -0.210 3.660 0.210 ;
        RECT  2.170 -0.210 2.290 0.500 ;
        RECT  1.490 -0.210 2.170 0.210 ;
        RECT  1.230 -0.210 1.490 0.260 ;
        RECT  0.680 -0.210 1.230 0.210 ;
        RECT  0.420 -0.210 0.680 0.230 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.115 2.310 12.320 2.730 ;
        RECT  11.945 1.480 12.115 2.730 ;
        RECT  11.395 2.310 11.945 2.730 ;
        RECT  11.225 1.740 11.395 2.730 ;
        RECT  10.570 2.310 11.225 2.730 ;
        RECT  10.140 1.960 10.570 2.730 ;
        RECT  8.090 2.310 10.140 2.730 ;
        RECT  7.920 1.910 8.090 2.730 ;
        RECT  7.280 2.310 7.920 2.730 ;
        RECT  7.110 1.910 7.280 2.730 ;
        RECT  6.315 2.310 7.110 2.730 ;
        RECT  6.055 2.190 6.315 2.730 ;
        RECT  4.785 2.310 6.055 2.730 ;
        RECT  4.615 2.260 4.785 2.730 ;
        RECT  4.295 2.310 4.615 2.730 ;
        RECT  4.125 2.260 4.295 2.730 ;
        RECT  2.625 2.310 4.125 2.730 ;
        RECT  2.365 2.290 2.625 2.730 ;
        RECT  1.595 2.310 2.365 2.730 ;
        RECT  1.335 2.260 1.595 2.730 ;
        RECT  0.530 2.310 1.335 2.730 ;
        RECT  0.360 2.265 0.530 2.730 ;
        RECT  0.000 2.310 0.360 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 12.320 2.520 ;
        LAYER M1 ;
        RECT  10.440 0.990 10.700 1.250 ;
        RECT  10.385 0.990 10.440 1.840 ;
        RECT  10.320 0.445 10.385 1.840 ;
        RECT  10.265 0.445 10.320 1.250 ;
        RECT  9.910 1.720 10.320 1.840 ;
        RECT  8.785 0.445 10.265 0.565 ;
        RECT  10.145 1.375 10.200 1.545 ;
        RECT  10.025 0.690 10.145 1.545 ;
        RECT  9.985 1.070 10.025 1.545 ;
        RECT  9.855 1.070 9.985 1.240 ;
        RECT  9.790 1.720 9.910 2.055 ;
        RECT  9.670 0.765 9.810 0.885 ;
        RECT  8.215 1.935 9.790 2.055 ;
        RECT  9.550 0.765 9.670 1.790 ;
        RECT  6.825 1.670 9.550 1.790 ;
        RECT  9.240 1.040 9.360 1.525 ;
        RECT  8.350 1.040 9.240 1.160 ;
        RECT  7.310 1.430 8.840 1.550 ;
        RECT  8.615 0.380 8.785 0.565 ;
        RECT  8.065 0.380 8.615 0.500 ;
        RECT  8.210 0.620 8.470 0.870 ;
        RECT  8.090 0.990 8.350 1.160 ;
        RECT  7.310 0.750 8.210 0.870 ;
        RECT  7.895 0.380 8.065 0.630 ;
        RECT  7.190 0.540 7.310 1.550 ;
        RECT  6.945 1.430 7.190 1.550 ;
        RECT  6.950 0.620 7.070 1.310 ;
        RECT  4.375 0.620 6.950 0.740 ;
        RECT  6.825 1.190 6.950 1.310 ;
        RECT  6.705 1.190 6.825 1.790 ;
        RECT  6.560 0.860 6.820 1.070 ;
        RECT  6.525 1.950 6.785 2.190 ;
        RECT  6.325 1.575 6.585 1.830 ;
        RECT  5.880 0.860 6.560 0.980 ;
        RECT  5.375 1.950 6.525 2.070 ;
        RECT  5.880 1.575 6.325 1.695 ;
        RECT  5.920 0.330 6.180 0.500 ;
        RECT  2.530 0.380 5.920 0.500 ;
        RECT  5.760 0.860 5.880 1.695 ;
        RECT  5.615 1.510 5.760 1.695 ;
        RECT  5.495 1.510 5.615 1.770 ;
        RECT  5.375 1.030 5.540 1.150 ;
        RECT  5.255 1.030 5.375 2.140 ;
        RECT  1.185 2.020 5.255 2.140 ;
        RECT  4.135 1.780 5.090 1.900 ;
        RECT  4.255 0.620 4.375 1.550 ;
        RECT  4.085 0.620 4.255 0.790 ;
        RECT  4.015 0.910 4.135 1.900 ;
        RECT  3.610 0.910 4.015 1.030 ;
        RECT  3.660 1.780 4.015 1.900 ;
        RECT  3.370 1.460 3.840 1.580 ;
        RECT  3.490 1.730 3.660 1.900 ;
        RECT  3.490 0.625 3.610 1.030 ;
        RECT  3.030 0.625 3.490 0.745 ;
        RECT  3.250 1.005 3.370 1.900 ;
        RECT  3.110 1.005 3.250 1.125 ;
        RECT  1.425 1.780 3.250 1.900 ;
        RECT  2.990 0.865 3.110 1.125 ;
        RECT  2.865 0.625 2.910 0.745 ;
        RECT  2.865 1.250 2.890 1.420 ;
        RECT  2.745 0.625 2.865 1.420 ;
        RECT  2.650 0.625 2.745 0.745 ;
        RECT  2.720 1.250 2.745 1.420 ;
        RECT  2.410 0.380 2.530 0.740 ;
        RECT  2.180 0.620 2.410 0.740 ;
        RECT  2.010 0.620 2.180 1.420 ;
        RECT  1.790 0.330 2.050 0.500 ;
        RECT  1.150 0.620 2.010 0.740 ;
        RECT  0.255 0.380 1.790 0.500 ;
        RECT  1.425 0.860 1.530 0.980 ;
        RECT  1.305 0.860 1.425 1.900 ;
        RECT  1.270 0.860 1.305 0.980 ;
        RECT  1.065 1.485 1.185 2.140 ;
        RECT  1.030 0.620 1.150 1.340 ;
        RECT  0.770 1.485 1.065 1.605 ;
        RECT  0.890 1.220 1.030 1.340 ;
        RECT  0.790 0.620 0.910 0.950 ;
        RECT  0.770 0.825 0.790 0.950 ;
        RECT  0.650 0.825 0.770 1.605 ;
        RECT  0.205 0.380 0.255 0.810 ;
        RECT  0.205 1.480 0.255 1.910 ;
        RECT  0.085 0.380 0.205 1.910 ;
    END
END SDFFSHQX8AD
MACRO SDFFSQX1AD
    CLASS CORE ;
    FOREIGN SDFFSQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.895 1.275 6.155 1.655 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.795 1.550 1.430 1.670 ;
        RECT  0.795 0.910 1.160 1.030 ;
        RECT  0.675 0.910 0.795 1.670 ;
        RECT  0.630 1.145 0.675 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.925 0.255 1.375 ;
        RECT  0.070 1.140 0.115 1.375 ;
        END
        AntennaGateArea 0.103 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.050 0.510 7.210 2.070 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 1.190 1.375 1.350 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.870 0.865 4.130 1.095 ;
        RECT  3.750 0.865 3.870 1.275 ;
        END
        AntennaGateArea 0.089 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.835 -0.210 7.280 0.210 ;
        RECT  6.665 -0.210 6.835 0.675 ;
        RECT  6.085 -0.210 6.665 0.210 ;
        RECT  5.915 -0.210 6.085 0.665 ;
        RECT  3.670 -0.210 5.915 0.210 ;
        RECT  3.410 -0.210 3.670 0.300 ;
        RECT  2.830 -0.210 3.410 0.210 ;
        RECT  2.570 -0.210 2.830 0.415 ;
        RECT  1.300 -0.210 2.570 0.210 ;
        RECT  1.040 -0.210 1.300 0.300 ;
        RECT  0.240 -0.210 1.040 0.210 ;
        RECT  0.120 -0.210 0.240 0.520 ;
        RECT  0.000 -0.210 0.120 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.825 2.310 7.280 2.730 ;
        RECT  6.565 2.015 6.825 2.730 ;
        RECT  5.840 2.310 6.565 2.730 ;
        RECT  5.670 2.055 5.840 2.730 ;
        RECT  4.800 2.310 5.670 2.730 ;
        RECT  4.540 2.020 4.800 2.730 ;
        RECT  4.010 2.310 4.540 2.730 ;
        RECT  3.750 1.965 4.010 2.730 ;
        RECT  2.685 2.310 3.750 2.730 ;
        RECT  2.565 1.995 2.685 2.730 ;
        RECT  1.245 2.310 2.565 2.730 ;
        RECT  1.075 2.050 1.245 2.730 ;
        RECT  0.240 2.310 1.075 2.730 ;
        RECT  0.120 1.880 0.240 2.730 ;
        RECT  0.000 2.310 0.120 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.280 2.520 ;
        LAYER M1 ;
        RECT  6.810 0.795 6.930 1.895 ;
        RECT  6.485 0.795 6.810 0.915 ;
        RECT  6.300 1.775 6.810 1.895 ;
        RECT  6.315 0.595 6.485 0.915 ;
        RECT  6.305 1.035 6.465 1.595 ;
        RECT  5.225 1.035 6.305 1.155 ;
        RECT  6.130 1.775 6.300 2.105 ;
        RECT  5.755 1.775 6.130 1.895 ;
        RECT  5.635 1.330 5.755 1.895 ;
        RECT  5.555 0.380 5.725 0.665 ;
        RECT  5.495 1.330 5.635 1.450 ;
        RECT  3.990 0.380 5.555 0.500 ;
        RECT  5.325 1.780 5.445 2.140 ;
        RECT  4.925 1.780 5.325 1.900 ;
        RECT  5.105 0.620 5.225 1.660 ;
        RECT  4.835 0.620 5.105 0.740 ;
        RECT  5.045 1.390 5.105 1.660 ;
        RECT  4.925 0.860 4.950 1.120 ;
        RECT  4.805 0.860 4.925 1.900 ;
        RECT  3.170 1.725 4.805 1.845 ;
        RECT  4.565 0.620 4.685 1.575 ;
        RECT  3.870 0.620 4.565 0.740 ;
        RECT  4.230 1.455 4.565 1.575 ;
        RECT  4.300 1.070 4.420 1.335 ;
        RECT  4.110 1.215 4.300 1.335 ;
        RECT  3.990 1.215 4.110 1.605 ;
        RECT  3.630 1.485 3.990 1.605 ;
        RECT  3.750 0.420 3.870 0.740 ;
        RECT  3.390 0.420 3.750 0.540 ;
        RECT  3.510 0.660 3.630 1.605 ;
        RECT  3.405 1.145 3.510 1.605 ;
        RECT  2.925 1.970 3.430 2.140 ;
        RECT  2.840 1.145 3.405 1.265 ;
        RECT  3.270 0.420 3.390 1.025 ;
        RECT  2.695 0.905 3.270 1.025 ;
        RECT  3.050 1.385 3.170 1.845 ;
        RECT  3.030 0.525 3.150 0.785 ;
        RECT  2.455 1.385 3.050 1.505 ;
        RECT  2.455 0.665 3.030 0.785 ;
        RECT  2.805 1.625 2.925 2.140 ;
        RECT  2.255 1.625 2.805 1.745 ;
        RECT  2.575 0.905 2.695 1.225 ;
        RECT  2.335 0.665 2.455 1.505 ;
        RECT  2.270 1.045 2.335 1.505 ;
        RECT  2.150 1.625 2.255 2.055 ;
        RECT  2.150 0.655 2.215 0.915 ;
        RECT  2.030 0.655 2.150 2.055 ;
        RECT  1.790 0.420 1.910 2.040 ;
        RECT  1.735 0.420 1.790 0.915 ;
        RECT  1.705 1.800 1.790 2.040 ;
        RECT  0.410 0.420 1.735 0.540 ;
        RECT  0.590 1.800 1.705 1.920 ;
        RECT  1.615 1.130 1.670 1.390 ;
        RECT  1.495 0.670 1.615 1.390 ;
        RECT  0.520 0.670 1.495 0.790 ;
        RECT  0.470 1.800 0.590 2.060 ;
        RECT  0.510 1.495 0.545 1.665 ;
        RECT  0.510 0.670 0.520 0.950 ;
        RECT  0.375 0.670 0.510 1.665 ;
    END
END SDFFSQX1AD
MACRO SDFFSQX2AD
    CLASS CORE ;
    FOREIGN SDFFSQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.890 1.275 6.155 1.655 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.795 1.550 1.430 1.670 ;
        RECT  0.795 0.910 1.160 1.030 ;
        RECT  0.675 0.910 0.795 1.670 ;
        RECT  0.630 1.145 0.675 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.925 0.255 1.375 ;
        RECT  0.070 1.140 0.115 1.375 ;
        END
        AntennaGateArea 0.103 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.050 0.380 7.210 1.985 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 1.190 1.375 1.350 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.870 0.865 4.130 1.095 ;
        RECT  3.750 0.865 3.870 1.275 ;
        END
        AntennaGateArea 0.088 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.835 -0.210 7.280 0.210 ;
        RECT  6.665 -0.210 6.835 0.575 ;
        RECT  6.085 -0.210 6.665 0.210 ;
        RECT  5.915 -0.210 6.085 0.655 ;
        RECT  3.670 -0.210 5.915 0.210 ;
        RECT  3.410 -0.210 3.670 0.300 ;
        RECT  2.830 -0.210 3.410 0.210 ;
        RECT  2.570 -0.210 2.830 0.415 ;
        RECT  1.300 -0.210 2.570 0.210 ;
        RECT  1.040 -0.210 1.300 0.300 ;
        RECT  0.230 -0.210 1.040 0.210 ;
        RECT  0.110 -0.210 0.230 0.520 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.825 2.310 7.280 2.730 ;
        RECT  6.565 2.015 6.825 2.730 ;
        RECT  5.840 2.310 6.565 2.730 ;
        RECT  5.670 2.055 5.840 2.730 ;
        RECT  4.800 2.310 5.670 2.730 ;
        RECT  4.540 2.020 4.800 2.730 ;
        RECT  4.010 2.310 4.540 2.730 ;
        RECT  3.750 1.965 4.010 2.730 ;
        RECT  2.685 2.310 3.750 2.730 ;
        RECT  2.565 1.995 2.685 2.730 ;
        RECT  1.245 2.310 2.565 2.730 ;
        RECT  1.075 2.050 1.245 2.730 ;
        RECT  0.240 2.310 1.075 2.730 ;
        RECT  0.120 1.880 0.240 2.730 ;
        RECT  0.000 2.310 0.120 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.280 2.520 ;
        LAYER M1 ;
        RECT  6.810 0.700 6.930 1.895 ;
        RECT  6.270 0.700 6.810 0.820 ;
        RECT  6.300 1.775 6.810 1.895 ;
        RECT  6.305 0.970 6.465 1.595 ;
        RECT  5.165 0.970 6.305 1.090 ;
        RECT  6.130 1.775 6.300 2.105 ;
        RECT  5.710 1.775 6.130 1.895 ;
        RECT  5.555 0.380 5.725 0.635 ;
        RECT  5.585 1.245 5.710 1.895 ;
        RECT  5.565 1.245 5.585 1.505 ;
        RECT  3.990 0.380 5.555 0.500 ;
        RECT  5.275 1.780 5.445 2.140 ;
        RECT  4.925 1.780 5.275 1.900 ;
        RECT  5.045 0.620 5.165 1.660 ;
        RECT  4.835 0.620 5.045 0.740 ;
        RECT  4.805 0.860 4.925 1.900 ;
        RECT  3.170 1.725 4.805 1.845 ;
        RECT  4.565 0.620 4.685 1.605 ;
        RECT  3.870 0.620 4.565 0.740 ;
        RECT  4.230 1.485 4.565 1.605 ;
        RECT  4.325 1.100 4.445 1.360 ;
        RECT  4.110 1.240 4.325 1.360 ;
        RECT  3.990 1.240 4.110 1.605 ;
        RECT  3.630 1.485 3.990 1.605 ;
        RECT  3.750 0.420 3.870 0.740 ;
        RECT  3.390 0.420 3.750 0.540 ;
        RECT  3.510 0.660 3.630 1.605 ;
        RECT  3.405 1.145 3.510 1.605 ;
        RECT  2.925 2.020 3.430 2.140 ;
        RECT  2.840 1.145 3.405 1.265 ;
        RECT  3.270 0.420 3.390 1.025 ;
        RECT  2.695 0.905 3.270 1.025 ;
        RECT  3.050 1.385 3.170 1.845 ;
        RECT  3.030 0.525 3.150 0.785 ;
        RECT  2.455 1.385 3.050 1.505 ;
        RECT  2.455 0.665 3.030 0.785 ;
        RECT  2.805 1.625 2.925 2.140 ;
        RECT  2.255 1.625 2.805 1.745 ;
        RECT  2.575 0.905 2.695 1.225 ;
        RECT  2.335 0.665 2.455 1.505 ;
        RECT  2.270 1.045 2.335 1.505 ;
        RECT  2.150 1.625 2.255 2.055 ;
        RECT  2.150 0.655 2.215 0.915 ;
        RECT  2.030 0.655 2.150 2.055 ;
        RECT  1.790 0.420 1.910 2.040 ;
        RECT  1.735 0.420 1.790 0.915 ;
        RECT  1.705 1.800 1.790 2.040 ;
        RECT  0.410 0.420 1.735 0.540 ;
        RECT  0.590 1.800 1.705 1.920 ;
        RECT  1.615 1.130 1.670 1.390 ;
        RECT  1.495 0.670 1.615 1.390 ;
        RECT  0.545 0.670 1.495 0.790 ;
        RECT  0.470 1.800 0.590 2.060 ;
        RECT  0.510 0.670 0.545 0.905 ;
        RECT  0.510 1.495 0.545 1.665 ;
        RECT  0.375 0.670 0.510 1.665 ;
    END
END SDFFSQX2AD
MACRO SDFFSQX4AD
    CLASS CORE ;
    FOREIGN SDFFSQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.895 1.275 6.155 1.655 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.795 1.550 1.430 1.670 ;
        RECT  0.795 0.910 1.160 1.030 ;
        RECT  0.675 0.910 0.795 1.670 ;
        RECT  0.630 1.145 0.675 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.925 0.255 1.375 ;
        RECT  0.070 1.140 0.115 1.375 ;
        END
        AntennaGateArea 0.103 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.070 0.425 7.210 1.985 ;
        RECT  6.945 0.425 7.070 0.855 ;
        RECT  6.970 1.465 7.070 1.985 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 1.190 1.375 1.350 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.870 0.865 4.130 1.095 ;
        RECT  3.750 0.865 3.870 1.280 ;
        END
        AntennaGateArea 0.088 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.450 -0.210 7.560 0.210 ;
        RECT  7.330 -0.210 7.450 0.840 ;
        RECT  6.755 -0.210 7.330 0.210 ;
        RECT  6.585 -0.210 6.755 0.485 ;
        RECT  6.085 -0.210 6.585 0.210 ;
        RECT  5.915 -0.210 6.085 0.655 ;
        RECT  3.670 -0.210 5.915 0.210 ;
        RECT  3.410 -0.210 3.670 0.300 ;
        RECT  2.830 -0.210 3.410 0.210 ;
        RECT  2.570 -0.210 2.830 0.415 ;
        RECT  1.300 -0.210 2.570 0.210 ;
        RECT  1.040 -0.210 1.300 0.300 ;
        RECT  0.240 -0.210 1.040 0.210 ;
        RECT  0.120 -0.210 0.240 0.520 ;
        RECT  0.000 -0.210 0.120 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.450 2.310 7.560 2.730 ;
        RECT  7.330 1.585 7.450 2.730 ;
        RECT  6.775 2.310 7.330 2.730 ;
        RECT  6.515 2.015 6.775 2.730 ;
        RECT  5.840 2.310 6.515 2.730 ;
        RECT  5.670 2.055 5.840 2.730 ;
        RECT  4.800 2.310 5.670 2.730 ;
        RECT  4.540 2.020 4.800 2.730 ;
        RECT  4.010 2.310 4.540 2.730 ;
        RECT  3.750 1.965 4.010 2.730 ;
        RECT  2.685 2.310 3.750 2.730 ;
        RECT  2.565 1.995 2.685 2.730 ;
        RECT  1.245 2.310 2.565 2.730 ;
        RECT  1.075 2.050 1.245 2.730 ;
        RECT  0.240 2.310 1.075 2.730 ;
        RECT  0.120 1.880 0.240 2.730 ;
        RECT  0.000 2.310 0.120 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  6.800 0.995 6.940 1.265 ;
        RECT  6.680 0.695 6.800 1.895 ;
        RECT  6.315 0.695 6.680 0.865 ;
        RECT  6.300 1.775 6.680 1.895 ;
        RECT  6.275 1.025 6.465 1.595 ;
        RECT  6.130 1.775 6.300 2.135 ;
        RECT  5.225 1.025 6.275 1.145 ;
        RECT  5.775 1.775 6.130 1.895 ;
        RECT  5.650 1.315 5.775 1.895 ;
        RECT  5.555 0.380 5.725 0.655 ;
        RECT  5.515 1.315 5.650 1.435 ;
        RECT  3.990 0.380 5.555 0.500 ;
        RECT  5.315 1.780 5.435 2.160 ;
        RECT  4.930 1.780 5.315 1.900 ;
        RECT  5.105 0.620 5.225 1.660 ;
        RECT  4.835 0.620 5.105 0.740 ;
        RECT  5.050 1.390 5.105 1.660 ;
        RECT  4.930 0.860 4.950 1.120 ;
        RECT  4.810 0.860 4.930 1.900 ;
        RECT  4.805 1.725 4.810 1.900 ;
        RECT  3.170 1.725 4.805 1.845 ;
        RECT  4.570 0.620 4.690 1.575 ;
        RECT  3.870 0.620 4.570 0.740 ;
        RECT  4.230 1.455 4.570 1.575 ;
        RECT  4.330 1.075 4.450 1.335 ;
        RECT  4.110 1.215 4.330 1.335 ;
        RECT  3.990 1.215 4.110 1.605 ;
        RECT  3.630 1.485 3.990 1.605 ;
        RECT  3.750 0.420 3.870 0.740 ;
        RECT  3.390 0.420 3.750 0.540 ;
        RECT  3.510 0.660 3.630 1.605 ;
        RECT  3.405 1.145 3.510 1.605 ;
        RECT  3.170 1.995 3.430 2.140 ;
        RECT  2.840 1.145 3.405 1.265 ;
        RECT  3.270 0.420 3.390 1.025 ;
        RECT  2.695 0.905 3.270 1.025 ;
        RECT  3.050 1.385 3.170 1.845 ;
        RECT  2.925 2.020 3.170 2.140 ;
        RECT  3.030 0.525 3.150 0.785 ;
        RECT  2.455 1.385 3.050 1.505 ;
        RECT  2.455 0.665 3.030 0.785 ;
        RECT  2.805 1.625 2.925 2.140 ;
        RECT  2.255 1.625 2.805 1.745 ;
        RECT  2.575 0.905 2.695 1.225 ;
        RECT  2.335 0.665 2.455 1.505 ;
        RECT  2.270 1.045 2.335 1.505 ;
        RECT  2.150 1.625 2.255 2.055 ;
        RECT  2.150 0.655 2.215 0.915 ;
        RECT  2.030 0.655 2.150 2.055 ;
        RECT  1.790 0.420 1.910 2.040 ;
        RECT  1.735 0.420 1.790 0.915 ;
        RECT  1.705 1.800 1.790 2.040 ;
        RECT  0.400 0.420 1.735 0.540 ;
        RECT  0.590 1.800 1.705 1.920 ;
        RECT  1.615 1.130 1.670 1.390 ;
        RECT  1.495 0.670 1.615 1.390 ;
        RECT  0.545 0.670 1.495 0.790 ;
        RECT  0.470 1.800 0.590 2.060 ;
        RECT  0.510 0.670 0.545 0.905 ;
        RECT  0.510 1.495 0.545 1.665 ;
        RECT  0.375 0.670 0.510 1.665 ;
    END
END SDFFSQX4AD
MACRO SDFFSQXLAD
    CLASS CORE ;
    FOREIGN SDFFSQXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.875 1.305 6.135 1.685 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.795 1.550 1.430 1.670 ;
        RECT  0.795 0.910 1.160 1.030 ;
        RECT  0.675 0.910 0.795 1.670 ;
        RECT  0.630 1.145 0.675 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.925 0.255 1.375 ;
        RECT  0.070 1.140 0.115 1.375 ;
        END
        AntennaGateArea 0.103 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.810 0.360 6.930 1.685 ;
        RECT  6.735 0.360 6.810 0.530 ;
        RECT  6.770 1.425 6.810 1.685 ;
        END
        AntennaDiffArea 0.142 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 1.190 1.375 1.350 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.870 0.865 4.130 1.095 ;
        RECT  3.750 0.865 3.870 1.275 ;
        END
        AntennaGateArea 0.087 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.545 -0.210 7.000 0.210 ;
        RECT  6.375 -0.210 6.545 0.530 ;
        RECT  6.065 -0.210 6.375 0.210 ;
        RECT  5.895 -0.210 6.065 0.665 ;
        RECT  3.690 -0.210 5.895 0.210 ;
        RECT  3.430 -0.210 3.690 0.300 ;
        RECT  2.830 -0.210 3.430 0.210 ;
        RECT  2.570 -0.210 2.830 0.415 ;
        RECT  1.300 -0.210 2.570 0.210 ;
        RECT  1.040 -0.210 1.300 0.300 ;
        RECT  0.240 -0.210 1.040 0.210 ;
        RECT  0.120 -0.210 0.240 0.520 ;
        RECT  0.000 -0.210 0.120 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.620 2.310 7.000 2.730 ;
        RECT  6.450 2.085 6.620 2.730 ;
        RECT  5.820 2.310 6.450 2.730 ;
        RECT  5.650 2.055 5.820 2.730 ;
        RECT  4.800 2.310 5.650 2.730 ;
        RECT  4.540 2.020 4.800 2.730 ;
        RECT  4.010 2.310 4.540 2.730 ;
        RECT  3.750 1.965 4.010 2.730 ;
        RECT  2.685 2.310 3.750 2.730 ;
        RECT  2.565 1.995 2.685 2.730 ;
        RECT  1.245 2.310 2.565 2.730 ;
        RECT  1.075 2.050 1.245 2.730 ;
        RECT  0.240 2.310 1.075 2.730 ;
        RECT  0.120 1.880 0.240 2.730 ;
        RECT  0.000 2.310 0.120 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.000 2.520 ;
        LAYER M1 ;
        RECT  6.630 1.005 6.665 1.265 ;
        RECT  6.510 0.725 6.630 1.935 ;
        RECT  6.270 0.725 6.510 0.845 ;
        RECT  6.230 1.815 6.510 1.935 ;
        RECT  5.225 1.005 6.390 1.125 ;
        RECT  6.060 1.815 6.230 1.985 ;
        RECT  5.685 1.815 6.060 1.935 ;
        RECT  5.535 0.380 5.705 0.765 ;
        RECT  5.565 1.245 5.685 1.935 ;
        RECT  3.990 0.380 5.535 0.500 ;
        RECT  5.300 1.780 5.425 2.140 ;
        RECT  4.925 1.780 5.300 1.900 ;
        RECT  5.105 0.620 5.225 1.650 ;
        RECT  4.835 0.620 5.105 0.740 ;
        RECT  5.045 1.390 5.105 1.650 ;
        RECT  4.925 0.860 4.950 1.120 ;
        RECT  4.805 0.860 4.925 1.900 ;
        RECT  3.170 1.725 4.805 1.845 ;
        RECT  4.565 0.620 4.685 1.575 ;
        RECT  3.870 0.620 4.565 0.740 ;
        RECT  4.230 1.455 4.565 1.575 ;
        RECT  4.300 1.070 4.420 1.335 ;
        RECT  4.110 1.215 4.300 1.335 ;
        RECT  3.990 1.215 4.110 1.605 ;
        RECT  3.630 1.485 3.990 1.605 ;
        RECT  3.750 0.420 3.870 0.740 ;
        RECT  3.390 0.420 3.750 0.540 ;
        RECT  3.510 0.660 3.630 1.605 ;
        RECT  3.405 1.145 3.510 1.605 ;
        RECT  2.925 1.970 3.430 2.140 ;
        RECT  2.840 1.145 3.405 1.265 ;
        RECT  3.270 0.420 3.390 1.025 ;
        RECT  2.695 0.905 3.270 1.025 ;
        RECT  3.050 1.385 3.170 1.845 ;
        RECT  3.030 0.525 3.150 0.785 ;
        RECT  2.455 1.385 3.050 1.505 ;
        RECT  2.455 0.665 3.030 0.785 ;
        RECT  2.805 1.625 2.925 2.140 ;
        RECT  2.255 1.625 2.805 1.745 ;
        RECT  2.575 0.905 2.695 1.225 ;
        RECT  2.335 0.665 2.455 1.505 ;
        RECT  2.270 1.045 2.335 1.505 ;
        RECT  2.150 1.625 2.255 2.055 ;
        RECT  2.150 0.655 2.215 0.915 ;
        RECT  2.030 0.655 2.150 2.055 ;
        RECT  1.790 0.420 1.910 2.040 ;
        RECT  1.735 0.420 1.790 0.915 ;
        RECT  1.705 1.800 1.790 2.040 ;
        RECT  0.410 0.420 1.735 0.540 ;
        RECT  0.590 1.800 1.705 1.920 ;
        RECT  1.615 1.130 1.670 1.390 ;
        RECT  1.495 0.670 1.615 1.390 ;
        RECT  0.520 0.670 1.495 0.790 ;
        RECT  0.470 1.800 0.590 2.060 ;
        RECT  0.510 1.495 0.545 1.665 ;
        RECT  0.510 0.670 0.520 0.950 ;
        RECT  0.375 0.670 0.510 1.665 ;
    END
END SDFFSQXLAD
MACRO SDFFSRHQX1AD
    CLASS CORE ;
    FOREIGN SDFFSRHQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.825 1.050 5.100 1.375 ;
        RECT  4.780 1.080 4.825 1.200 ;
        END
        AntennaGateArea 0.109 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.775 1.030 4.175 1.330 ;
        END
        AntennaGateArea 0.05 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 1.280 3.370 1.660 ;
        RECT  1.890 1.540 3.250 1.660 ;
        RECT  1.520 1.145 1.890 1.660 ;
        END
        AntennaGateArea 0.098 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.215 1.020 9.335 1.280 ;
        RECT  8.050 1.080 9.215 1.200 ;
        RECT  7.910 1.080 8.050 1.375 ;
        END
        AntennaGateArea 0.101 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.370 1.145 11.410 1.375 ;
        RECT  11.250 0.615 11.370 1.890 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 0.865 2.810 1.130 ;
        END
        AntennaGateArea 0.053 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.930 0.490 1.375 ;
        END
        AntennaGateArea 0.12 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.060 -0.210 11.480 0.210 ;
        RECT  10.800 -0.210 11.060 0.310 ;
        RECT  9.835 -0.210 10.800 0.210 ;
        RECT  9.575 -0.210 9.835 0.310 ;
        RECT  8.075 -0.210 9.575 0.210 ;
        RECT  7.815 -0.210 8.075 0.300 ;
        RECT  6.845 -0.210 7.815 0.210 ;
        RECT  6.585 -0.210 6.845 0.300 ;
        RECT  5.010 -0.210 6.585 0.210 ;
        RECT  4.750 -0.210 5.010 0.300 ;
        RECT  4.200 -0.210 4.750 0.210 ;
        RECT  3.940 -0.210 4.200 0.300 ;
        RECT  2.510 -0.210 3.940 0.210 ;
        RECT  2.250 -0.210 2.510 0.260 ;
        RECT  1.315 -0.210 2.250 0.210 ;
        RECT  1.055 -0.210 1.315 0.260 ;
        RECT  0.680 -0.210 1.055 0.210 ;
        RECT  0.420 -0.210 0.680 0.260 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.050 2.310 11.480 2.730 ;
        RECT  10.790 2.010 11.050 2.730 ;
        RECT  9.595 2.310 10.790 2.730 ;
        RECT  9.335 2.220 9.595 2.730 ;
        RECT  7.905 2.310 9.335 2.730 ;
        RECT  7.645 2.260 7.905 2.730 ;
        RECT  7.245 2.310 7.645 2.730 ;
        RECT  6.985 2.260 7.245 2.730 ;
        RECT  6.365 2.310 6.985 2.730 ;
        RECT  6.105 2.260 6.365 2.730 ;
        RECT  4.805 2.310 6.105 2.730 ;
        RECT  4.545 2.260 4.805 2.730 ;
        RECT  2.710 2.310 4.545 2.730 ;
        RECT  2.450 2.260 2.710 2.730 ;
        RECT  1.950 2.310 2.450 2.730 ;
        RECT  1.690 2.260 1.950 2.730 ;
        RECT  0.570 2.310 1.690 2.730 ;
        RECT  0.350 1.880 0.570 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.480 2.520 ;
        LAYER M1 ;
        RECT  11.015 1.000 11.120 1.260 ;
        RECT  10.895 0.430 11.015 1.885 ;
        RECT  8.945 0.430 10.895 0.550 ;
        RECT  10.740 1.000 10.895 1.260 ;
        RECT  10.525 1.765 10.895 1.885 ;
        RECT  10.600 0.695 10.695 0.815 ;
        RECT  10.455 0.695 10.600 1.590 ;
        RECT  10.265 1.765 10.525 2.025 ;
        RECT  9.815 0.695 10.455 0.815 ;
        RECT  10.195 1.160 10.315 1.645 ;
        RECT  8.775 1.905 10.265 2.025 ;
        RECT  9.575 1.160 10.195 1.280 ;
        RECT  9.160 1.400 10.075 1.575 ;
        RECT  9.695 0.695 9.815 1.040 ;
        RECT  9.455 0.780 9.575 1.280 ;
        RECT  8.565 0.780 9.455 0.900 ;
        RECT  8.945 1.400 9.160 1.785 ;
        RECT  8.685 0.430 8.945 0.660 ;
        RECT  8.560 1.665 8.945 1.785 ;
        RECT  8.290 1.425 8.655 1.545 ;
        RECT  6.825 2.020 8.655 2.140 ;
        RECT  8.445 0.420 8.565 0.900 ;
        RECT  8.410 1.665 8.560 1.860 ;
        RECT  6.195 0.420 8.445 0.540 ;
        RECT  7.035 1.740 8.410 1.860 ;
        RECT  7.275 0.680 8.325 0.805 ;
        RECT  8.170 1.425 8.290 1.620 ;
        RECT  7.275 1.500 8.170 1.620 ;
        RECT  7.155 0.680 7.275 1.620 ;
        RECT  6.915 0.660 7.035 1.860 ;
        RECT  4.655 0.660 6.915 0.780 ;
        RECT  6.565 2.020 6.825 2.185 ;
        RECT  6.660 0.900 6.735 1.160 ;
        RECT  6.660 1.715 6.705 1.835 ;
        RECT  6.490 0.900 6.660 1.835 ;
        RECT  5.515 2.020 6.565 2.140 ;
        RECT  5.700 0.900 6.490 1.020 ;
        RECT  5.755 1.715 6.490 1.835 ;
        RECT  5.935 0.380 6.195 0.540 ;
        RECT  3.710 0.420 5.935 0.540 ;
        RECT  5.635 1.540 5.755 1.835 ;
        RECT  5.395 0.990 5.515 2.140 ;
        RECT  5.305 0.990 5.395 1.250 ;
        RECT  1.150 2.020 5.395 2.140 ;
        RECT  4.415 1.740 5.275 1.860 ;
        RECT  4.535 0.660 4.655 1.590 ;
        RECT  4.295 0.660 4.415 1.860 ;
        RECT  3.470 0.660 4.295 0.780 ;
        RECT  3.730 1.740 4.295 1.860 ;
        RECT  3.610 1.450 4.110 1.570 ;
        RECT  3.590 0.380 3.710 0.540 ;
        RECT  3.490 0.900 3.610 1.900 ;
        RECT  2.225 0.380 3.590 0.500 ;
        RECT  3.180 0.900 3.490 1.160 ;
        RECT  1.390 1.780 3.490 1.900 ;
        RECT  3.210 0.620 3.470 0.780 ;
        RECT  3.060 1.300 3.100 1.420 ;
        RECT  2.930 0.620 3.060 1.420 ;
        RECT  2.770 0.620 2.930 0.740 ;
        RECT  2.840 1.300 2.930 1.420 ;
        RECT  2.225 1.300 2.430 1.420 ;
        RECT  2.105 0.380 2.225 1.420 ;
        RECT  1.140 0.620 2.105 0.740 ;
        RECT  1.600 0.330 1.860 0.500 ;
        RECT  1.390 0.860 1.790 0.980 ;
        RECT  0.230 0.380 1.600 0.500 ;
        RECT  1.270 0.860 1.390 1.900 ;
        RECT  1.030 1.460 1.150 2.140 ;
        RECT  1.020 0.620 1.140 1.270 ;
        RECT  0.730 1.460 1.030 1.580 ;
        RECT  0.850 1.095 1.020 1.270 ;
        RECT  0.730 0.660 0.900 0.920 ;
        RECT  0.610 0.660 0.730 1.580 ;
        RECT  0.110 0.380 0.230 1.600 ;
    END
END SDFFSRHQX1AD
MACRO SDFFSRHQX2AD
    CLASS CORE ;
    FOREIGN SDFFSRHQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.825 1.050 5.100 1.375 ;
        RECT  4.780 1.080 4.825 1.200 ;
        END
        AntennaGateArea 0.131 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.775 1.030 4.175 1.330 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 1.280 3.370 1.620 ;
        RECT  1.935 1.500 3.250 1.620 ;
        RECT  1.750 1.470 1.935 1.620 ;
        RECT  1.510 1.215 1.750 1.620 ;
        END
        AntennaGateArea 0.096 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.215 1.020 9.335 1.280 ;
        RECT  8.050 1.080 9.215 1.200 ;
        RECT  7.910 1.080 8.050 1.375 ;
        END
        AntennaGateArea 0.131 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.370 1.145 11.410 1.375 ;
        RECT  11.250 0.370 11.370 1.990 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 0.865 2.840 1.130 ;
        END
        AntennaGateArea 0.081 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.930 0.490 1.375 ;
        END
        AntennaGateArea 0.116 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.010 -0.210 11.480 0.210 ;
        RECT  10.750 -0.210 11.010 0.310 ;
        RECT  9.835 -0.210 10.750 0.210 ;
        RECT  9.575 -0.210 9.835 0.310 ;
        RECT  8.075 -0.210 9.575 0.210 ;
        RECT  7.815 -0.210 8.075 0.300 ;
        RECT  6.845 -0.210 7.815 0.210 ;
        RECT  6.585 -0.210 6.845 0.300 ;
        RECT  5.015 -0.210 6.585 0.210 ;
        RECT  4.755 -0.210 5.015 0.300 ;
        RECT  4.205 -0.210 4.755 0.210 ;
        RECT  3.945 -0.210 4.205 0.300 ;
        RECT  2.470 -0.210 3.945 0.210 ;
        RECT  2.350 -0.210 2.470 0.390 ;
        RECT  1.315 -0.210 2.350 0.210 ;
        RECT  1.055 -0.210 1.315 0.300 ;
        RECT  0.680 -0.210 1.055 0.210 ;
        RECT  0.420 -0.210 0.680 0.300 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.050 2.310 11.480 2.730 ;
        RECT  10.790 2.010 11.050 2.730 ;
        RECT  9.685 2.310 10.790 2.730 ;
        RECT  9.425 2.220 9.685 2.730 ;
        RECT  7.995 2.310 9.425 2.730 ;
        RECT  7.735 2.225 7.995 2.730 ;
        RECT  7.245 2.310 7.735 2.730 ;
        RECT  6.985 2.225 7.245 2.730 ;
        RECT  6.455 2.310 6.985 2.730 ;
        RECT  6.195 2.225 6.455 2.730 ;
        RECT  4.795 2.310 6.195 2.730 ;
        RECT  4.535 2.225 4.795 2.730 ;
        RECT  2.850 2.310 4.535 2.730 ;
        RECT  2.590 2.225 2.850 2.730 ;
        RECT  1.950 2.310 2.590 2.730 ;
        RECT  1.690 2.225 1.950 2.730 ;
        RECT  0.570 2.310 1.690 2.730 ;
        RECT  0.350 1.880 0.570 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.480 2.520 ;
        LAYER M1 ;
        RECT  11.015 1.000 11.120 1.260 ;
        RECT  10.895 0.430 11.015 1.885 ;
        RECT  8.945 0.430 10.895 0.550 ;
        RECT  10.740 1.000 10.895 1.260 ;
        RECT  10.525 1.765 10.895 1.885 ;
        RECT  10.620 0.695 10.650 0.905 ;
        RECT  10.455 0.695 10.620 1.590 ;
        RECT  10.265 1.765 10.525 2.045 ;
        RECT  9.815 0.695 10.455 0.815 ;
        RECT  10.185 1.160 10.305 1.645 ;
        RECT  8.775 1.925 10.265 2.045 ;
        RECT  9.575 1.160 10.185 1.280 ;
        RECT  9.160 1.400 10.065 1.575 ;
        RECT  9.695 0.695 9.815 1.040 ;
        RECT  9.455 0.780 9.575 1.280 ;
        RECT  8.565 0.780 9.455 0.900 ;
        RECT  8.945 1.400 9.160 1.805 ;
        RECT  8.685 0.430 8.945 0.660 ;
        RECT  8.560 1.675 8.945 1.805 ;
        RECT  8.290 1.435 8.655 1.555 ;
        RECT  8.445 0.420 8.565 0.900 ;
        RECT  8.410 1.675 8.560 1.865 ;
        RECT  8.205 1.985 8.465 2.190 ;
        RECT  6.195 0.420 8.445 0.540 ;
        RECT  7.035 1.745 8.410 1.865 ;
        RECT  7.300 0.680 8.325 0.805 ;
        RECT  8.170 1.435 8.290 1.615 ;
        RECT  6.825 1.985 8.205 2.105 ;
        RECT  7.300 1.495 8.170 1.615 ;
        RECT  7.155 0.680 7.300 1.615 ;
        RECT  6.915 0.660 7.035 1.865 ;
        RECT  4.655 0.660 6.915 0.780 ;
        RECT  6.565 1.985 6.825 2.170 ;
        RECT  6.660 0.900 6.735 1.160 ;
        RECT  6.660 1.690 6.705 1.810 ;
        RECT  6.490 0.900 6.660 1.835 ;
        RECT  5.515 1.985 6.565 2.105 ;
        RECT  5.705 0.900 6.490 1.020 ;
        RECT  6.445 1.690 6.490 1.835 ;
        RECT  5.755 1.715 6.445 1.835 ;
        RECT  5.935 0.380 6.195 0.540 ;
        RECT  3.710 0.420 5.935 0.540 ;
        RECT  5.635 1.540 5.755 1.835 ;
        RECT  5.395 0.990 5.515 2.105 ;
        RECT  5.305 0.990 5.395 1.250 ;
        RECT  1.150 1.985 5.395 2.105 ;
        RECT  4.415 1.740 5.275 1.860 ;
        RECT  4.535 0.660 4.655 1.590 ;
        RECT  4.295 0.660 4.415 1.860 ;
        RECT  3.470 0.660 4.295 0.780 ;
        RECT  3.730 1.740 4.295 1.860 ;
        RECT  3.610 1.450 4.110 1.570 ;
        RECT  3.590 0.380 3.710 0.540 ;
        RECT  3.490 0.900 3.610 1.860 ;
        RECT  2.710 0.380 3.590 0.500 ;
        RECT  3.210 0.900 3.490 1.160 ;
        RECT  1.390 1.740 3.490 1.860 ;
        RECT  3.210 0.620 3.470 0.780 ;
        RECT  3.090 1.260 3.130 1.380 ;
        RECT  2.960 0.620 3.090 1.380 ;
        RECT  2.830 0.620 2.960 0.740 ;
        RECT  2.870 1.260 2.960 1.380 ;
        RECT  2.590 0.380 2.710 0.705 ;
        RECT  2.225 0.585 2.590 0.705 ;
        RECT  2.225 1.260 2.460 1.380 ;
        RECT  2.105 0.585 2.225 1.380 ;
        RECT  1.935 0.585 2.105 0.780 ;
        RECT  1.140 0.660 1.935 0.780 ;
        RECT  1.645 0.335 1.815 0.540 ;
        RECT  1.390 0.900 1.800 1.020 ;
        RECT  0.230 0.420 1.645 0.540 ;
        RECT  1.270 0.900 1.390 1.860 ;
        RECT  1.030 1.460 1.150 2.105 ;
        RECT  1.020 0.660 1.140 1.260 ;
        RECT  0.730 1.460 1.030 1.580 ;
        RECT  0.850 1.090 1.020 1.260 ;
        RECT  0.730 0.660 0.900 0.920 ;
        RECT  0.610 0.660 0.730 1.580 ;
        RECT  0.110 0.420 0.230 1.600 ;
    END
END SDFFSRHQX2AD
MACRO SDFFSRHQX4AD
    CLASS CORE ;
    FOREIGN SDFFSRHQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.720 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.825 1.050 5.100 1.375 ;
        RECT  4.780 1.080 4.825 1.200 ;
        END
        AntennaGateArea 0.159 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 1.030 4.175 1.330 ;
        END
        AntennaGateArea 0.072 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 1.280 3.370 1.620 ;
        RECT  1.935 1.500 3.250 1.620 ;
        RECT  1.750 1.470 1.935 1.620 ;
        RECT  1.510 1.215 1.750 1.620 ;
        END
        AntennaGateArea 0.12 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.270 1.025 11.415 1.330 ;
        RECT  10.050 1.190 11.270 1.330 ;
        RECT  9.885 1.190 10.050 1.380 ;
        RECT  9.200 1.260 9.885 1.380 ;
        END
        AntennaGateArea 0.215 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.230 0.355 13.370 2.040 ;
        RECT  13.130 0.355 13.230 0.875 ;
        RECT  13.130 1.520 13.230 2.040 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 0.865 2.840 1.130 ;
        END
        AntennaGateArea 0.14 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.930 0.490 1.375 ;
        END
        AntennaGateArea 0.172 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.610 -0.210 13.720 0.210 ;
        RECT  13.490 -0.210 13.610 0.875 ;
        RECT  12.760 -0.210 13.490 0.210 ;
        RECT  12.590 -0.210 12.760 0.260 ;
        RECT  11.860 -0.210 12.590 0.210 ;
        RECT  11.690 -0.210 11.860 0.260 ;
        RECT  9.105 -0.210 11.690 0.210 ;
        RECT  8.845 -0.210 9.105 0.630 ;
        RECT  7.895 -0.210 8.845 0.210 ;
        RECT  7.635 -0.210 7.895 0.300 ;
        RECT  6.955 -0.210 7.635 0.210 ;
        RECT  6.695 -0.210 6.955 0.300 ;
        RECT  5.015 -0.210 6.695 0.210 ;
        RECT  4.755 -0.210 5.015 0.300 ;
        RECT  4.215 -0.210 4.755 0.210 ;
        RECT  3.955 -0.210 4.215 0.300 ;
        RECT  2.470 -0.210 3.955 0.210 ;
        RECT  2.350 -0.210 2.470 0.390 ;
        RECT  1.315 -0.210 2.350 0.210 ;
        RECT  1.055 -0.210 1.315 0.300 ;
        RECT  0.680 -0.210 1.055 0.210 ;
        RECT  0.420 -0.210 0.680 0.300 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.610 2.310 13.720 2.730 ;
        RECT  13.490 1.590 13.610 2.730 ;
        RECT  12.940 2.310 13.490 2.730 ;
        RECT  12.680 2.010 12.940 2.730 ;
        RECT  11.520 2.310 12.680 2.730 ;
        RECT  11.260 2.210 11.520 2.730 ;
        RECT  8.860 2.310 11.260 2.730 ;
        RECT  8.430 2.260 8.860 2.730 ;
        RECT  7.785 2.310 8.430 2.730 ;
        RECT  7.615 2.260 7.785 2.730 ;
        RECT  6.525 2.310 7.615 2.730 ;
        RECT  6.265 1.890 6.525 2.730 ;
        RECT  4.945 2.310 6.265 2.730 ;
        RECT  4.425 2.220 4.945 2.730 ;
        RECT  2.740 2.310 4.425 2.730 ;
        RECT  2.480 2.220 2.740 2.730 ;
        RECT  1.950 2.310 2.480 2.730 ;
        RECT  1.690 2.220 1.950 2.730 ;
        RECT  0.570 2.310 1.690 2.730 ;
        RECT  0.350 2.050 0.570 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 13.720 2.520 ;
        LAYER M1 ;
        RECT  12.900 1.000 13.065 1.260 ;
        RECT  12.780 0.380 12.900 1.890 ;
        RECT  10.005 0.380 12.780 0.500 ;
        RECT  12.685 1.000 12.780 1.260 ;
        RECT  12.440 1.770 12.780 1.890 ;
        RECT  12.565 0.710 12.590 0.905 ;
        RECT  12.445 0.710 12.565 1.590 ;
        RECT  12.420 0.710 12.445 0.905 ;
        RECT  12.270 1.770 12.440 2.085 ;
        RECT  11.895 0.710 12.420 0.835 ;
        RECT  12.120 1.090 12.290 1.635 ;
        RECT  11.110 1.965 12.270 2.085 ;
        RECT  11.655 1.090 12.120 1.210 ;
        RECT  11.845 1.360 11.965 1.620 ;
        RECT  11.775 0.710 11.895 0.970 ;
        RECT  10.870 1.460 11.845 1.580 ;
        RECT  11.535 0.660 11.655 1.210 ;
        RECT  9.415 0.660 11.535 0.780 ;
        RECT  10.990 1.965 11.110 2.140 ;
        RECT  9.960 2.020 10.990 2.140 ;
        RECT  10.750 1.460 10.870 1.900 ;
        RECT  9.090 1.780 10.750 1.900 ;
        RECT  9.785 0.900 10.645 1.020 ;
        RECT  9.690 1.540 10.610 1.660 ;
        RECT  9.585 0.900 9.785 1.110 ;
        RECT  9.430 1.500 9.690 1.660 ;
        RECT  7.415 2.020 9.670 2.140 ;
        RECT  8.425 0.990 9.585 1.110 ;
        RECT  8.425 1.500 9.430 1.620 ;
        RECT  9.295 0.660 9.415 0.870 ;
        RECT  8.665 0.750 9.295 0.870 ;
        RECT  8.970 1.740 9.090 1.900 ;
        RECT  7.380 1.740 8.970 1.860 ;
        RECT  8.545 0.420 8.665 0.870 ;
        RECT  7.345 0.420 8.545 0.540 ;
        RECT  8.305 0.660 8.425 1.620 ;
        RECT  7.970 1.385 8.305 1.620 ;
        RECT  8.045 0.660 8.165 1.260 ;
        RECT  4.655 0.660 8.045 0.780 ;
        RECT  7.380 1.140 8.045 1.260 ;
        RECT  7.500 1.385 7.970 1.505 ;
        RECT  7.035 0.900 7.925 1.020 ;
        RECT  7.155 2.020 7.415 2.185 ;
        RECT  7.260 1.140 7.380 1.860 ;
        RECT  7.085 0.340 7.345 0.540 ;
        RECT  6.765 2.020 7.155 2.140 ;
        RECT  7.035 1.635 7.140 1.895 ;
        RECT  3.835 0.420 7.085 0.540 ;
        RECT  6.915 0.900 7.035 1.895 ;
        RECT  5.695 0.900 6.915 1.020 ;
        RECT  5.755 1.405 6.915 1.525 ;
        RECT  6.645 1.645 6.765 2.140 ;
        RECT  5.995 1.645 6.645 1.765 ;
        RECT  5.515 1.140 6.470 1.260 ;
        RECT  5.875 1.645 5.995 2.125 ;
        RECT  5.515 2.005 5.875 2.125 ;
        RECT  5.635 1.405 5.755 1.885 ;
        RECT  5.395 0.990 5.515 2.125 ;
        RECT  5.305 0.990 5.395 1.260 ;
        RECT  1.150 1.980 5.395 2.100 ;
        RECT  4.415 1.740 5.275 1.860 ;
        RECT  4.535 0.660 4.655 1.590 ;
        RECT  4.295 0.660 4.415 1.860 ;
        RECT  3.500 0.660 4.295 0.780 ;
        RECT  3.730 1.740 4.295 1.860 ;
        RECT  3.610 1.450 4.110 1.570 ;
        RECT  3.715 0.380 3.835 0.540 ;
        RECT  2.710 0.380 3.715 0.500 ;
        RECT  3.490 0.900 3.610 1.860 ;
        RECT  3.240 0.620 3.500 0.780 ;
        RECT  3.230 0.900 3.490 1.160 ;
        RECT  1.390 1.740 3.490 1.860 ;
        RECT  3.090 1.260 3.130 1.380 ;
        RECT  2.960 0.620 3.090 1.380 ;
        RECT  2.830 0.620 2.960 0.740 ;
        RECT  2.870 1.260 2.960 1.380 ;
        RECT  2.590 0.380 2.710 0.705 ;
        RECT  2.225 0.585 2.590 0.705 ;
        RECT  2.225 1.260 2.460 1.380 ;
        RECT  2.105 0.585 2.225 1.380 ;
        RECT  1.935 0.585 2.105 0.780 ;
        RECT  1.140 0.660 1.935 0.780 ;
        RECT  1.815 0.360 1.860 0.480 ;
        RECT  1.600 0.360 1.815 0.540 ;
        RECT  1.390 0.900 1.800 1.020 ;
        RECT  0.230 0.420 1.600 0.540 ;
        RECT  1.270 0.900 1.390 1.860 ;
        RECT  1.030 1.460 1.150 2.100 ;
        RECT  1.020 0.660 1.140 1.235 ;
        RECT  0.730 1.460 1.030 1.580 ;
        RECT  0.850 1.060 1.020 1.235 ;
        RECT  0.730 0.660 0.900 0.920 ;
        RECT  0.610 0.660 0.730 1.580 ;
        RECT  0.110 0.420 0.230 1.600 ;
    END
END SDFFSRHQX4AD
MACRO SDFFSRHQX8AD
    CLASS CORE ;
    FOREIGN SDFFSRHQX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.825 1.035 5.100 1.375 ;
        END
        AntennaGateArea 0.184 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 1.030 4.175 1.330 ;
        END
        AntennaGateArea 0.108 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 1.280 3.370 1.620 ;
        RECT  1.935 1.500 3.250 1.620 ;
        RECT  1.690 1.190 1.935 1.620 ;
        END
        AntennaGateArea 0.173 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.295 1.070 11.415 1.330 ;
        RECT  10.050 1.190 11.295 1.330 ;
        RECT  9.885 1.190 10.050 1.380 ;
        RECT  9.085 1.260 9.885 1.380 ;
        END
        AntennaGateArea 0.25 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.935 0.355 14.105 2.125 ;
        RECT  13.440 1.005 13.935 1.515 ;
        RECT  13.240 0.400 13.440 2.125 ;
        RECT  13.215 0.400 13.240 0.830 ;
        RECT  13.215 1.435 13.240 2.125 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.545 0.865 2.830 1.130 ;
        END
        AntennaGateArea 0.16 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.930 0.490 1.375 ;
        END
        AntennaGateArea 0.266 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.440 -0.210 14.560 0.210 ;
        RECT  14.320 -0.210 14.440 0.875 ;
        RECT  13.720 -0.210 14.320 0.210 ;
        RECT  13.600 -0.210 13.720 0.875 ;
        RECT  13.000 -0.210 13.600 0.210 ;
        RECT  12.740 -0.210 13.000 0.350 ;
        RECT  11.955 -0.210 12.740 0.210 ;
        RECT  11.695 -0.210 11.955 0.300 ;
        RECT  9.170 -0.210 11.695 0.210 ;
        RECT  8.910 -0.210 9.170 0.630 ;
        RECT  7.895 -0.210 8.910 0.210 ;
        RECT  7.635 -0.210 7.895 0.300 ;
        RECT  6.955 -0.210 7.635 0.210 ;
        RECT  6.695 -0.210 6.955 0.300 ;
        RECT  5.015 -0.210 6.695 0.210 ;
        RECT  4.755 -0.210 5.015 0.300 ;
        RECT  4.220 -0.210 4.755 0.210 ;
        RECT  3.960 -0.210 4.220 0.260 ;
        RECT  2.730 -0.210 3.960 0.210 ;
        RECT  2.470 -0.210 2.730 0.255 ;
        RECT  1.425 -0.210 2.470 0.210 ;
        RECT  1.165 -0.210 1.425 0.300 ;
        RECT  0.680 -0.210 1.165 0.210 ;
        RECT  0.420 -0.210 0.680 0.300 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.465 2.310 14.560 2.730 ;
        RECT  14.295 1.435 14.465 2.730 ;
        RECT  13.780 2.310 14.295 2.730 ;
        RECT  13.580 1.700 13.780 2.730 ;
        RECT  13.070 2.310 13.580 2.730 ;
        RECT  12.810 2.040 13.070 2.730 ;
        RECT  11.625 2.310 12.810 2.730 ;
        RECT  11.365 2.230 11.625 2.730 ;
        RECT  8.610 2.310 11.365 2.730 ;
        RECT  8.350 2.220 8.610 2.730 ;
        RECT  7.830 2.310 8.350 2.730 ;
        RECT  7.570 2.220 7.830 2.730 ;
        RECT  6.585 2.310 7.570 2.730 ;
        RECT  6.325 1.890 6.585 2.730 ;
        RECT  5.010 2.310 6.325 2.730 ;
        RECT  4.490 2.260 5.010 2.730 ;
        RECT  2.705 2.310 4.490 2.730 ;
        RECT  2.535 2.265 2.705 2.730 ;
        RECT  1.985 2.310 2.535 2.730 ;
        RECT  1.725 2.220 1.985 2.730 ;
        RECT  0.570 2.310 1.725 2.730 ;
        RECT  0.350 2.050 0.570 2.730 ;
        RECT  0.000 2.310 0.350 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 14.560 2.520 ;
        LAYER M1 ;
        RECT  12.940 1.045 13.120 1.215 ;
        RECT  12.940 1.800 12.945 1.920 ;
        RECT  12.790 0.470 12.940 1.920 ;
        RECT  12.370 0.470 12.790 0.590 ;
        RECT  12.690 1.045 12.790 1.215 ;
        RECT  12.440 1.800 12.790 1.920 ;
        RECT  12.570 0.735 12.640 0.905 ;
        RECT  12.410 0.735 12.570 1.590 ;
        RECT  12.225 1.800 12.440 2.085 ;
        RECT  11.895 0.785 12.410 0.905 ;
        RECT  12.200 0.355 12.370 0.590 ;
        RECT  12.120 1.180 12.290 1.680 ;
        RECT  11.235 1.905 12.225 2.085 ;
        RECT  12.030 0.420 12.200 0.590 ;
        RECT  11.655 1.180 12.120 1.300 ;
        RECT  11.025 0.420 12.030 0.540 ;
        RECT  11.845 1.420 11.965 1.680 ;
        RECT  11.775 0.785 11.895 1.060 ;
        RECT  10.975 1.460 11.845 1.580 ;
        RECT  11.535 0.830 11.655 1.300 ;
        RECT  11.030 0.830 11.535 0.950 ;
        RECT  11.115 1.905 11.235 2.140 ;
        RECT  9.945 2.020 11.115 2.140 ;
        RECT  10.910 0.660 11.030 0.950 ;
        RECT  10.765 0.380 11.025 0.540 ;
        RECT  10.855 1.460 10.975 1.900 ;
        RECT  10.075 0.660 10.910 0.780 ;
        RECT  9.090 1.780 10.855 1.900 ;
        RECT  10.005 0.380 10.765 0.500 ;
        RECT  9.760 0.900 10.645 1.020 ;
        RECT  9.690 1.540 10.565 1.660 ;
        RECT  9.815 0.620 10.075 0.780 ;
        RECT  9.440 0.660 9.815 0.780 ;
        RECT  9.600 0.900 9.760 1.110 ;
        RECT  9.430 1.500 9.690 1.660 ;
        RECT  8.850 2.020 9.655 2.140 ;
        RECT  8.965 0.990 9.600 1.110 ;
        RECT  9.300 0.660 9.440 0.870 ;
        RECT  8.965 1.500 9.430 1.620 ;
        RECT  8.665 0.750 9.300 0.870 ;
        RECT  8.970 1.740 9.090 1.900 ;
        RECT  8.725 1.740 8.970 1.860 ;
        RECT  8.845 0.990 8.965 1.620 ;
        RECT  8.730 1.980 8.850 2.140 ;
        RECT  8.425 0.990 8.845 1.110 ;
        RECT  7.415 1.980 8.730 2.100 ;
        RECT  8.605 1.300 8.725 1.860 ;
        RECT  8.545 0.420 8.665 0.870 ;
        RECT  7.380 1.740 8.605 1.860 ;
        RECT  7.345 0.420 8.545 0.540 ;
        RECT  8.305 0.660 8.425 1.620 ;
        RECT  7.970 1.385 8.305 1.620 ;
        RECT  8.045 0.660 8.165 1.260 ;
        RECT  4.655 0.660 8.045 0.780 ;
        RECT  7.380 1.140 8.045 1.260 ;
        RECT  7.500 1.385 7.970 1.505 ;
        RECT  7.140 0.900 7.925 1.020 ;
        RECT  7.275 1.980 7.415 2.185 ;
        RECT  7.260 1.140 7.380 1.860 ;
        RECT  7.085 0.330 7.345 0.540 ;
        RECT  7.155 2.020 7.275 2.185 ;
        RECT  6.885 2.020 7.155 2.140 ;
        RECT  7.020 0.900 7.140 1.895 ;
        RECT  4.665 0.420 7.085 0.540 ;
        RECT  5.695 0.900 7.020 1.020 ;
        RECT  5.885 1.405 7.020 1.525 ;
        RECT  6.765 1.645 6.885 2.140 ;
        RECT  6.150 1.645 6.765 1.765 ;
        RECT  5.645 1.140 6.470 1.260 ;
        RECT  6.030 1.645 6.150 2.140 ;
        RECT  5.645 2.020 6.030 2.140 ;
        RECT  5.765 1.405 5.885 1.860 ;
        RECT  5.525 1.140 5.645 2.140 ;
        RECT  5.425 1.140 5.525 1.260 ;
        RECT  3.555 2.020 5.525 2.140 ;
        RECT  5.305 0.990 5.425 1.260 ;
        RECT  4.415 1.780 5.375 1.900 ;
        RECT  4.545 0.380 4.665 0.540 ;
        RECT  4.535 0.660 4.655 1.570 ;
        RECT  2.380 0.380 4.545 0.500 ;
        RECT  4.295 0.620 4.415 1.900 ;
        RECT  3.280 0.620 4.295 0.740 ;
        RECT  3.730 1.780 4.295 1.900 ;
        RECT  3.610 1.450 4.110 1.570 ;
        RECT  3.490 0.900 3.610 1.860 ;
        RECT  3.305 1.980 3.555 2.140 ;
        RECT  3.215 0.900 3.490 1.160 ;
        RECT  1.570 1.740 3.490 1.860 ;
        RECT  1.205 1.980 3.305 2.100 ;
        RECT  3.090 0.620 3.160 0.740 ;
        RECT  3.090 1.260 3.130 1.380 ;
        RECT  2.950 0.620 3.090 1.380 ;
        RECT  2.900 0.620 2.950 0.740 ;
        RECT  2.870 1.260 2.950 1.380 ;
        RECT  2.380 1.260 2.450 1.380 ;
        RECT  2.260 0.380 2.380 1.380 ;
        RECT  2.110 0.380 2.260 0.780 ;
        RECT  2.190 1.260 2.260 1.380 ;
        RECT  1.330 0.660 2.110 0.780 ;
        RECT  1.680 0.370 1.850 0.540 ;
        RECT  1.570 0.900 1.810 1.020 ;
        RECT  0.230 0.420 1.680 0.540 ;
        RECT  1.450 0.900 1.570 1.860 ;
        RECT  1.345 1.740 1.450 1.860 ;
        RECT  1.210 0.660 1.330 1.235 ;
        RECT  1.025 1.060 1.210 1.235 ;
        RECT  1.050 1.460 1.205 2.100 ;
        RECT  0.900 0.660 1.060 0.830 ;
        RECT  0.900 1.460 1.050 1.580 ;
        RECT  0.780 0.660 0.900 1.580 ;
        RECT  0.110 0.380 0.230 1.940 ;
    END
END SDFFSRHQX8AD
MACRO SDFFSRX1AD
    CLASS CORE ;
    FOREIGN SDFFSRX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.585 0.955 7.820 1.395 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 0.950 1.460 1.810 ;
        RECT  1.145 0.950 1.340 1.330 ;
        RECT  1.000 0.950 1.145 1.210 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.050 0.485 1.220 ;
        RECT  0.070 1.050 0.210 1.375 ;
        END
        AntennaGateArea 0.103 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.980 4.410 1.440 ;
        END
        AntennaGateArea 0.048 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.690 1.360 8.890 1.655 ;
        RECT  8.525 0.680 8.690 1.655 ;
        END
        AntennaDiffArea 0.207 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.290 0.615 9.450 1.890 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.865 1.460 1.190 1.760 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.985 1.025 4.130 1.540 ;
        END
        AntennaGateArea 0.083 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.075 -0.210 9.520 0.210 ;
        RECT  8.905 -0.210 9.075 0.825 ;
        RECT  8.005 -0.210 8.905 0.210 ;
        RECT  7.835 -0.210 8.005 0.525 ;
        RECT  4.310 -0.210 7.835 0.210 ;
        RECT  4.050 -0.210 4.310 0.300 ;
        RECT  2.995 -0.210 4.050 0.210 ;
        RECT  2.825 -0.210 2.995 0.650 ;
        RECT  1.360 -0.210 2.825 0.210 ;
        RECT  1.100 -0.210 1.360 0.310 ;
        RECT  0.275 -0.210 1.100 0.210 ;
        RECT  0.105 -0.210 0.275 0.905 ;
        RECT  0.000 -0.210 0.105 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.100 2.310 9.520 2.730 ;
        RECT  8.840 2.015 9.100 2.730 ;
        RECT  8.365 2.310 8.840 2.730 ;
        RECT  8.105 2.015 8.365 2.730 ;
        RECT  6.420 2.310 8.105 2.730 ;
        RECT  6.160 2.210 6.420 2.730 ;
        RECT  4.880 2.310 6.160 2.730 ;
        RECT  4.620 2.040 4.880 2.730 ;
        RECT  4.220 2.310 4.620 2.730 ;
        RECT  3.960 2.075 4.220 2.730 ;
        RECT  2.960 2.310 3.960 2.730 ;
        RECT  2.840 1.995 2.960 2.730 ;
        RECT  1.315 2.310 2.840 2.730 ;
        RECT  1.145 2.170 1.315 2.730 ;
        RECT  0.275 2.310 1.145 2.730 ;
        RECT  0.110 1.495 0.275 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.520 2.520 ;
        LAYER M1 ;
        RECT  9.050 1.020 9.170 1.895 ;
        RECT  8.405 1.775 9.050 1.895 ;
        RECT  8.285 0.355 8.405 1.895 ;
        RECT  8.195 0.355 8.285 0.525 ;
        RECT  7.235 1.515 8.285 1.690 ;
        RECT  8.005 0.670 8.125 1.365 ;
        RECT  6.520 0.670 8.005 0.790 ;
        RECT  5.515 0.380 7.690 0.500 ;
        RECT  7.270 1.855 7.530 2.090 ;
        RECT  5.020 1.970 7.270 2.090 ;
        RECT  6.835 0.960 7.005 1.850 ;
        RECT  6.640 0.960 6.835 1.115 ;
        RECT  4.890 1.730 6.835 1.850 ;
        RECT  6.520 1.480 6.695 1.600 ;
        RECT  6.400 0.670 6.520 1.600 ;
        RECT  6.160 0.890 6.280 1.600 ;
        RECT  6.030 0.890 6.160 1.010 ;
        RECT  5.460 1.480 6.160 1.600 ;
        RECT  5.035 1.200 6.040 1.320 ;
        RECT  5.770 0.830 6.030 1.010 ;
        RECT  5.275 0.890 5.770 1.010 ;
        RECT  5.395 0.380 5.515 0.770 ;
        RECT  5.155 0.420 5.275 1.010 ;
        RECT  3.625 0.420 5.155 0.540 ;
        RECT  4.915 0.660 5.035 1.320 ;
        RECT  3.890 0.660 4.915 0.780 ;
        RECT  4.770 1.730 4.890 1.920 ;
        RECT  4.715 0.900 4.790 1.020 ;
        RECT  4.245 1.800 4.770 1.920 ;
        RECT  4.650 0.900 4.715 1.430 ;
        RECT  4.530 0.900 4.650 1.680 ;
        RECT  4.370 1.560 4.530 1.680 ;
        RECT  4.125 1.730 4.245 1.920 ;
        RECT  3.440 1.730 4.125 1.850 ;
        RECT  3.865 0.660 3.890 0.920 ;
        RECT  3.745 0.660 3.865 1.610 ;
        RECT  3.575 1.255 3.745 1.610 ;
        RECT  3.505 0.420 3.625 1.135 ;
        RECT  3.200 2.020 3.600 2.140 ;
        RECT  2.970 1.255 3.575 1.375 ;
        RECT  2.790 1.015 3.505 1.135 ;
        RECT  3.320 1.515 3.440 1.850 ;
        RECT  3.215 0.715 3.385 0.890 ;
        RECT  2.540 1.515 3.320 1.635 ;
        RECT  2.540 0.770 3.215 0.890 ;
        RECT  3.080 1.755 3.200 2.140 ;
        RECT  2.305 1.755 3.080 1.875 ;
        RECT  2.670 1.015 2.790 1.285 ;
        RECT  2.420 0.770 2.540 1.635 ;
        RECT  2.370 1.255 2.420 1.635 ;
        RECT  2.250 1.755 2.305 2.075 ;
        RECT  2.250 0.670 2.300 0.930 ;
        RECT  2.130 0.670 2.250 2.075 ;
        RECT  1.940 0.810 2.010 2.050 ;
        RECT  1.890 0.430 1.940 2.050 ;
        RECT  1.820 0.430 1.890 0.930 ;
        RECT  0.685 1.930 1.890 2.050 ;
        RECT  0.730 0.430 1.820 0.550 ;
        RECT  1.700 1.140 1.770 1.660 ;
        RECT  1.650 0.710 1.700 1.660 ;
        RECT  1.580 0.710 1.650 1.330 ;
        RECT  0.730 0.710 1.580 0.830 ;
        RECT  0.470 0.375 0.730 0.550 ;
        RECT  0.605 0.710 0.730 1.555 ;
        RECT  0.515 1.930 0.685 2.100 ;
        RECT  0.465 0.735 0.605 0.905 ;
        RECT  0.465 1.385 0.605 1.555 ;
    END
END SDFFSRX1AD
MACRO SDFFSRX2AD
    CLASS CORE ;
    FOREIGN SDFFSRX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.865 0.955 8.100 1.395 ;
        END
        AntennaGateArea 0.101 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 0.950 1.460 1.810 ;
        RECT  1.145 0.950 1.340 1.330 ;
        RECT  1.000 0.950 1.145 1.210 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.050 0.485 1.220 ;
        RECT  0.070 1.050 0.210 1.375 ;
        END
        AntennaGateArea 0.103 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.880 4.410 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.970 1.360 9.170 1.655 ;
        RECT  8.805 0.415 8.970 1.655 ;
        END
        AntennaDiffArea 0.373 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.690 0.615 9.730 1.985 ;
        RECT  9.570 0.415 9.690 1.985 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.865 1.460 1.190 1.760 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.965 0.990 4.130 1.540 ;
        END
        AntennaGateArea 0.096 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.355 -0.210 9.800 0.210 ;
        RECT  9.185 -0.210 9.355 0.810 ;
        RECT  8.285 -0.210 9.185 0.210 ;
        RECT  8.115 -0.210 8.285 0.525 ;
        RECT  4.285 -0.210 8.115 0.210 ;
        RECT  4.025 -0.210 4.285 0.260 ;
        RECT  2.985 -0.210 4.025 0.210 ;
        RECT  2.815 -0.210 2.985 0.650 ;
        RECT  1.360 -0.210 2.815 0.210 ;
        RECT  1.100 -0.210 1.360 0.300 ;
        RECT  0.275 -0.210 1.100 0.210 ;
        RECT  0.105 -0.210 0.275 0.905 ;
        RECT  0.000 -0.210 0.105 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.380 2.310 9.800 2.730 ;
        RECT  9.120 2.035 9.380 2.730 ;
        RECT  8.645 2.310 9.120 2.730 ;
        RECT  8.385 2.015 8.645 2.730 ;
        RECT  6.815 2.310 8.385 2.730 ;
        RECT  6.555 2.260 6.815 2.730 ;
        RECT  4.805 2.310 6.555 2.730 ;
        RECT  4.545 2.220 4.805 2.730 ;
        RECT  4.220 2.310 4.545 2.730 ;
        RECT  3.960 2.220 4.220 2.730 ;
        RECT  2.960 2.310 3.960 2.730 ;
        RECT  2.840 1.995 2.960 2.730 ;
        RECT  1.315 2.310 2.840 2.730 ;
        RECT  1.145 2.170 1.315 2.730 ;
        RECT  0.275 2.310 1.145 2.730 ;
        RECT  0.110 1.495 0.275 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.800 2.520 ;
        LAYER M1 ;
        RECT  9.330 1.020 9.450 1.895 ;
        RECT  8.685 1.775 9.330 1.895 ;
        RECT  8.565 0.355 8.685 1.895 ;
        RECT  8.475 0.355 8.565 0.525 ;
        RECT  7.500 1.515 8.565 1.690 ;
        RECT  8.285 0.670 8.405 1.380 ;
        RECT  6.575 0.670 8.285 0.790 ;
        RECT  5.510 0.380 7.970 0.500 ;
        RECT  7.695 1.855 7.835 1.975 ;
        RECT  7.575 1.855 7.695 2.140 ;
        RECT  5.595 2.020 7.575 2.140 ;
        RECT  7.195 0.960 7.315 1.900 ;
        RECT  6.915 0.960 7.195 1.080 ;
        RECT  5.835 1.780 7.195 1.900 ;
        RECT  6.575 1.480 6.995 1.600 ;
        RECT  6.455 0.670 6.575 1.600 ;
        RECT  6.215 0.890 6.335 1.520 ;
        RECT  6.200 0.890 6.215 1.010 ;
        RECT  6.075 1.400 6.215 1.520 ;
        RECT  5.680 0.830 6.200 1.010 ;
        RECT  5.030 1.160 6.095 1.280 ;
        RECT  5.955 1.400 6.075 1.660 ;
        RECT  5.715 1.440 5.835 1.900 ;
        RECT  4.935 1.440 5.715 1.560 ;
        RECT  5.270 0.890 5.680 1.010 ;
        RECT  5.475 1.690 5.595 2.140 ;
        RECT  5.390 0.380 5.510 0.770 ;
        RECT  5.075 1.690 5.475 1.810 ;
        RECT  5.235 1.930 5.355 2.190 ;
        RECT  5.150 0.380 5.270 1.010 ;
        RECT  3.200 1.980 5.235 2.100 ;
        RECT  3.605 0.380 5.150 0.500 ;
        RECT  4.910 0.620 5.030 1.280 ;
        RECT  4.815 1.440 4.935 1.860 ;
        RECT  3.845 0.620 4.910 0.740 ;
        RECT  3.440 1.740 4.815 1.860 ;
        RECT  4.740 0.860 4.790 0.980 ;
        RECT  4.650 0.860 4.740 1.310 ;
        RECT  4.530 0.860 4.650 1.620 ;
        RECT  4.345 1.500 4.530 1.620 ;
        RECT  3.725 0.620 3.845 1.610 ;
        RECT  3.575 1.255 3.725 1.610 ;
        RECT  3.485 0.380 3.605 1.135 ;
        RECT  2.970 1.255 3.575 1.375 ;
        RECT  2.790 1.015 3.485 1.135 ;
        RECT  3.320 1.515 3.440 1.860 ;
        RECT  3.195 0.715 3.365 0.890 ;
        RECT  2.540 1.515 3.320 1.635 ;
        RECT  3.080 1.755 3.200 2.100 ;
        RECT  2.540 0.770 3.195 0.890 ;
        RECT  2.305 1.755 3.080 1.875 ;
        RECT  2.670 1.015 2.790 1.285 ;
        RECT  2.420 0.770 2.540 1.635 ;
        RECT  2.370 1.255 2.420 1.635 ;
        RECT  2.250 1.755 2.305 2.075 ;
        RECT  2.250 0.670 2.300 0.930 ;
        RECT  2.180 0.670 2.250 2.075 ;
        RECT  2.130 0.735 2.180 2.075 ;
        RECT  1.940 0.810 2.010 2.050 ;
        RECT  1.890 0.420 1.940 2.050 ;
        RECT  1.820 0.420 1.890 0.930 ;
        RECT  0.685 1.930 1.890 2.050 ;
        RECT  0.470 0.420 1.820 0.540 ;
        RECT  1.700 1.140 1.770 1.660 ;
        RECT  1.650 0.710 1.700 1.660 ;
        RECT  1.580 0.710 1.650 1.330 ;
        RECT  0.730 0.710 1.580 0.830 ;
        RECT  0.605 0.710 0.730 1.555 ;
        RECT  0.515 1.930 0.685 2.100 ;
        RECT  0.465 0.735 0.605 0.905 ;
        RECT  0.465 1.385 0.605 1.555 ;
    END
END SDFFSRX2AD
MACRO SDFFSRX4AD
    CLASS CORE ;
    FOREIGN SDFFSRX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.115 1.190 9.540 1.420 ;
        END
        AntennaGateArea 0.15 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 0.950 1.460 1.810 ;
        RECT  1.145 0.950 1.340 1.330 ;
        RECT  1.000 0.950 1.145 1.210 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.050 0.485 1.220 ;
        RECT  0.070 1.050 0.210 1.375 ;
        END
        AntennaGateArea 0.106 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.880 4.410 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.430 0.415 10.570 1.655 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.330 1.005 11.410 1.515 ;
        RECT  11.170 0.415 11.330 1.985 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.865 1.460 1.190 1.760 ;
        END
        AntennaGateArea 0.065 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.965 0.990 4.130 1.540 ;
        END
        AntennaGateArea 0.119 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.675 -0.210 11.760 0.210 ;
        RECT  11.505 -0.210 11.675 0.810 ;
        RECT  10.955 -0.210 11.505 0.210 ;
        RECT  10.785 -0.210 10.955 0.810 ;
        RECT  10.235 -0.210 10.785 0.210 ;
        RECT  10.065 -0.210 10.235 0.415 ;
        RECT  9.255 -0.210 10.065 0.210 ;
        RECT  9.085 -0.210 9.255 0.575 ;
        RECT  4.285 -0.210 9.085 0.210 ;
        RECT  4.025 -0.210 4.285 0.260 ;
        RECT  2.985 -0.210 4.025 0.210 ;
        RECT  2.815 -0.210 2.985 0.650 ;
        RECT  1.360 -0.210 2.815 0.210 ;
        RECT  1.100 -0.210 1.360 0.300 ;
        RECT  0.275 -0.210 1.100 0.210 ;
        RECT  0.105 -0.210 0.275 0.905 ;
        RECT  0.000 -0.210 0.105 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.675 2.310 11.760 2.730 ;
        RECT  11.505 1.780 11.675 2.730 ;
        RECT  11.000 2.310 11.505 2.730 ;
        RECT  10.740 2.035 11.000 2.730 ;
        RECT  10.280 2.310 10.740 2.730 ;
        RECT  10.020 2.015 10.280 2.730 ;
        RECT  8.340 2.310 10.020 2.730 ;
        RECT  8.080 2.260 8.340 2.730 ;
        RECT  5.650 2.310 8.080 2.730 ;
        RECT  5.480 2.220 5.650 2.730 ;
        RECT  4.855 2.310 5.480 2.730 ;
        RECT  4.595 2.220 4.855 2.730 ;
        RECT  4.220 2.310 4.595 2.730 ;
        RECT  3.960 2.220 4.220 2.730 ;
        RECT  2.960 2.310 3.960 2.730 ;
        RECT  2.840 1.995 2.960 2.730 ;
        RECT  1.315 2.310 2.840 2.730 ;
        RECT  1.145 2.170 1.315 2.730 ;
        RECT  0.275 2.310 1.145 2.730 ;
        RECT  0.110 1.495 0.275 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.760 2.520 ;
        LAYER M1 ;
        RECT  10.930 1.020 11.050 1.895 ;
        RECT  10.310 1.775 10.930 1.895 ;
        RECT  10.190 0.710 10.310 1.895 ;
        RECT  9.680 0.710 10.190 0.830 ;
        RECT  9.065 1.540 10.190 1.725 ;
        RECT  9.885 0.950 10.005 1.260 ;
        RECT  8.500 0.950 9.885 1.070 ;
        RECT  9.520 0.370 9.660 0.490 ;
        RECT  9.400 0.370 9.520 0.830 ;
        RECT  8.895 0.710 9.400 0.830 ;
        RECT  9.230 1.890 9.400 2.010 ;
        RECT  9.110 1.890 9.230 2.140 ;
        RECT  6.880 2.020 9.110 2.140 ;
        RECT  8.775 0.530 8.895 0.830 ;
        RECT  8.760 1.510 8.880 1.860 ;
        RECT  8.725 0.530 8.775 0.765 ;
        RECT  8.230 1.740 8.760 1.860 ;
        RECT  8.620 0.530 8.725 0.650 ;
        RECT  8.500 1.500 8.640 1.620 ;
        RECT  8.500 0.380 8.620 0.650 ;
        RECT  6.070 0.380 8.500 0.500 ;
        RECT  8.380 0.770 8.500 1.620 ;
        RECT  8.310 0.770 8.380 0.890 ;
        RECT  8.050 0.620 8.310 0.890 ;
        RECT  8.110 1.010 8.230 1.860 ;
        RECT  7.950 1.010 8.110 1.130 ;
        RECT  6.505 1.740 8.110 1.860 ;
        RECT  7.830 0.770 8.050 0.890 ;
        RECT  7.710 0.620 7.830 1.620 ;
        RECT  6.950 0.620 7.710 0.740 ;
        RECT  7.340 1.500 7.710 1.620 ;
        RECT  7.220 0.860 7.590 0.980 ;
        RECT  7.100 0.860 7.220 1.620 ;
        RECT  6.430 0.860 7.100 0.980 ;
        RECT  6.960 1.500 7.100 1.620 ;
        RECT  6.860 1.100 6.980 1.360 ;
        RECT  6.620 1.980 6.880 2.140 ;
        RECT  5.155 1.160 6.860 1.280 ;
        RECT  6.130 2.020 6.620 2.140 ;
        RECT  6.385 1.440 6.505 1.860 ;
        RECT  6.170 0.810 6.430 0.980 ;
        RECT  4.895 1.440 6.385 1.560 ;
        RECT  5.640 0.860 6.170 0.980 ;
        RECT  6.010 1.690 6.130 2.140 ;
        RECT  5.950 0.380 6.070 0.740 ;
        RECT  5.055 1.690 6.010 1.810 ;
        RECT  5.810 0.620 5.950 0.740 ;
        RECT  5.770 1.930 5.890 2.190 ;
        RECT  3.200 1.980 5.770 2.100 ;
        RECT  5.520 0.380 5.640 0.980 ;
        RECT  3.605 0.380 5.520 0.500 ;
        RECT  5.035 0.620 5.155 1.280 ;
        RECT  3.845 0.620 5.035 0.740 ;
        RECT  4.775 1.440 4.895 1.860 ;
        RECT  4.740 0.860 4.790 0.980 ;
        RECT  3.450 1.740 4.775 1.860 ;
        RECT  4.650 0.860 4.740 1.310 ;
        RECT  4.530 0.860 4.650 1.620 ;
        RECT  4.345 1.500 4.530 1.620 ;
        RECT  3.725 0.620 3.845 1.610 ;
        RECT  3.575 1.255 3.725 1.610 ;
        RECT  3.485 0.380 3.605 1.135 ;
        RECT  2.970 1.255 3.575 1.375 ;
        RECT  2.790 1.015 3.485 1.135 ;
        RECT  3.330 1.515 3.450 1.860 ;
        RECT  3.195 0.715 3.365 0.890 ;
        RECT  2.540 1.515 3.330 1.635 ;
        RECT  3.080 1.755 3.200 2.100 ;
        RECT  2.540 0.770 3.195 0.890 ;
        RECT  2.305 1.755 3.080 1.875 ;
        RECT  2.670 1.015 2.790 1.285 ;
        RECT  2.420 0.770 2.540 1.635 ;
        RECT  2.370 1.255 2.420 1.635 ;
        RECT  2.250 1.755 2.305 2.075 ;
        RECT  2.250 0.670 2.300 0.930 ;
        RECT  2.130 0.670 2.250 2.075 ;
        RECT  1.940 0.810 2.010 2.050 ;
        RECT  1.890 0.420 1.940 2.050 ;
        RECT  1.820 0.420 1.890 0.930 ;
        RECT  0.685 1.930 1.890 2.050 ;
        RECT  0.470 0.420 1.820 0.540 ;
        RECT  1.700 1.140 1.770 1.660 ;
        RECT  1.650 0.710 1.700 1.660 ;
        RECT  1.580 0.710 1.650 1.330 ;
        RECT  0.730 0.710 1.580 0.830 ;
        RECT  0.605 0.710 0.730 1.555 ;
        RECT  0.515 1.930 0.685 2.100 ;
        RECT  0.465 0.735 0.605 0.905 ;
        RECT  0.465 1.385 0.605 1.555 ;
    END
END SDFFSRX4AD
MACRO SDFFSRXLAD
    CLASS CORE ;
    FOREIGN SDFFSRXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.585 0.955 7.820 1.395 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 0.950 1.460 1.810 ;
        RECT  1.145 0.950 1.340 1.330 ;
        RECT  1.000 0.950 1.145 1.210 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.050 0.485 1.220 ;
        RECT  0.070 1.050 0.210 1.375 ;
        END
        AntennaGateArea 0.103 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.980 4.410 1.440 ;
        END
        AntennaGateArea 0.048 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.410 1.360 8.610 1.655 ;
        RECT  8.245 0.680 8.410 1.655 ;
        END
        AntennaDiffArea 0.143 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.010 0.675 9.170 1.670 ;
        END
        AntennaDiffArea 0.143 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.865 1.460 1.190 1.760 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.985 1.025 4.130 1.540 ;
        END
        AntennaGateArea 0.083 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.860 -0.210 9.240 0.210 ;
        RECT  8.600 -0.210 8.860 0.320 ;
        RECT  8.005 -0.210 8.600 0.210 ;
        RECT  7.835 -0.210 8.005 0.525 ;
        RECT  4.310 -0.210 7.835 0.210 ;
        RECT  4.050 -0.210 4.310 0.300 ;
        RECT  2.995 -0.210 4.050 0.210 ;
        RECT  2.825 -0.210 2.995 0.650 ;
        RECT  1.360 -0.210 2.825 0.210 ;
        RECT  1.100 -0.210 1.360 0.310 ;
        RECT  0.275 -0.210 1.100 0.210 ;
        RECT  0.105 -0.210 0.275 0.905 ;
        RECT  0.000 -0.210 0.105 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.820 2.310 9.240 2.730 ;
        RECT  8.560 2.015 8.820 2.730 ;
        RECT  8.345 2.310 8.560 2.730 ;
        RECT  8.085 2.015 8.345 2.730 ;
        RECT  6.420 2.310 8.085 2.730 ;
        RECT  6.160 2.210 6.420 2.730 ;
        RECT  4.880 2.310 6.160 2.730 ;
        RECT  4.620 2.040 4.880 2.730 ;
        RECT  4.220 2.310 4.620 2.730 ;
        RECT  3.960 2.075 4.220 2.730 ;
        RECT  2.960 2.310 3.960 2.730 ;
        RECT  2.840 1.995 2.960 2.730 ;
        RECT  1.315 2.310 2.840 2.730 ;
        RECT  1.145 2.170 1.315 2.730 ;
        RECT  0.275 2.310 1.145 2.730 ;
        RECT  0.110 1.495 0.275 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.240 2.520 ;
        LAYER M1 ;
        RECT  8.770 0.440 8.890 1.895 ;
        RECT  8.365 0.440 8.770 0.560 ;
        RECT  7.915 1.775 8.770 1.895 ;
        RECT  8.235 0.355 8.365 0.560 ;
        RECT  8.195 0.355 8.235 0.525 ;
        RECT  8.005 0.670 8.125 1.365 ;
        RECT  6.520 0.670 8.005 0.790 ;
        RECT  7.795 1.565 7.915 2.135 ;
        RECT  7.405 1.565 7.795 1.685 ;
        RECT  5.515 0.380 7.690 0.500 ;
        RECT  7.270 1.855 7.530 2.090 ;
        RECT  7.235 1.515 7.405 1.685 ;
        RECT  5.020 1.970 7.270 2.090 ;
        RECT  6.835 0.960 7.005 1.850 ;
        RECT  6.640 0.960 6.835 1.115 ;
        RECT  4.890 1.730 6.835 1.850 ;
        RECT  6.520 1.480 6.695 1.600 ;
        RECT  6.400 0.670 6.520 1.600 ;
        RECT  6.160 0.890 6.280 1.600 ;
        RECT  6.030 0.890 6.160 1.010 ;
        RECT  5.460 1.480 6.160 1.600 ;
        RECT  5.035 1.200 6.040 1.320 ;
        RECT  5.770 0.830 6.030 1.010 ;
        RECT  5.275 0.890 5.770 1.010 ;
        RECT  5.395 0.380 5.515 0.770 ;
        RECT  5.155 0.420 5.275 1.010 ;
        RECT  3.625 0.420 5.155 0.540 ;
        RECT  4.915 0.660 5.035 1.320 ;
        RECT  3.890 0.660 4.915 0.780 ;
        RECT  4.770 1.730 4.890 1.920 ;
        RECT  4.715 0.900 4.790 1.020 ;
        RECT  4.245 1.800 4.770 1.920 ;
        RECT  4.650 0.900 4.715 1.430 ;
        RECT  4.530 0.900 4.650 1.680 ;
        RECT  4.370 1.560 4.530 1.680 ;
        RECT  4.125 1.730 4.245 1.920 ;
        RECT  3.440 1.730 4.125 1.850 ;
        RECT  3.865 0.660 3.890 0.920 ;
        RECT  3.745 0.660 3.865 1.610 ;
        RECT  3.575 1.255 3.745 1.610 ;
        RECT  3.505 0.420 3.625 1.135 ;
        RECT  3.200 2.020 3.600 2.140 ;
        RECT  2.970 1.255 3.575 1.375 ;
        RECT  2.790 1.015 3.505 1.135 ;
        RECT  3.320 1.515 3.440 1.850 ;
        RECT  3.215 0.715 3.385 0.890 ;
        RECT  2.540 1.515 3.320 1.635 ;
        RECT  2.540 0.770 3.215 0.890 ;
        RECT  3.080 1.755 3.200 2.140 ;
        RECT  2.305 1.755 3.080 1.875 ;
        RECT  2.670 1.015 2.790 1.285 ;
        RECT  2.420 0.770 2.540 1.635 ;
        RECT  2.370 1.255 2.420 1.635 ;
        RECT  2.250 1.755 2.305 2.075 ;
        RECT  2.250 0.670 2.300 0.930 ;
        RECT  2.130 0.670 2.250 2.075 ;
        RECT  1.940 0.810 2.010 2.050 ;
        RECT  1.890 0.430 1.940 2.050 ;
        RECT  1.820 0.430 1.890 0.930 ;
        RECT  0.685 1.930 1.890 2.050 ;
        RECT  0.730 0.430 1.820 0.550 ;
        RECT  1.700 1.140 1.770 1.660 ;
        RECT  1.650 0.710 1.700 1.660 ;
        RECT  1.580 0.710 1.650 1.330 ;
        RECT  0.730 0.710 1.580 0.830 ;
        RECT  0.470 0.375 0.730 0.550 ;
        RECT  0.605 0.710 0.730 1.555 ;
        RECT  0.515 1.930 0.685 2.100 ;
        RECT  0.465 0.735 0.605 0.905 ;
        RECT  0.465 1.385 0.605 1.555 ;
    END
END SDFFSRXLAD
MACRO SDFFSX1AD
    CLASS CORE ;
    FOREIGN SDFFSX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.910 1.100 6.090 1.620 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 1.560 1.430 1.680 ;
        RECT  0.995 0.930 1.160 1.070 ;
        RECT  0.875 0.930 0.995 1.680 ;
        RECT  0.630 1.145 0.875 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.265 1.280 ;
        RECT  0.070 1.020 0.210 1.655 ;
        END
        AntennaGateArea 0.103 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.670 0.690 6.780 0.950 ;
        RECT  6.670 1.330 6.780 1.590 ;
        RECT  6.510 0.690 6.670 1.590 ;
        END
        AntennaDiffArea 0.168 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.350 0.640 7.490 1.895 ;
        RECT  7.320 0.640 7.350 0.900 ;
        RECT  7.320 1.375 7.350 1.895 ;
        END
        AntennaDiffArea 0.203 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 1.190 1.415 1.430 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.925 0.910 4.175 1.090 ;
        RECT  3.805 0.910 3.925 1.275 ;
        END
        AntennaGateArea 0.089 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.265 -0.210 7.560 0.210 ;
        RECT  7.145 -0.210 7.265 0.420 ;
        RECT  6.240 -0.210 7.145 0.210 ;
        RECT  5.980 -0.210 6.240 0.310 ;
        RECT  4.005 -0.210 5.980 0.210 ;
        RECT  3.835 -0.210 4.005 0.370 ;
        RECT  2.710 -0.210 3.835 0.210 ;
        RECT  2.450 -0.210 2.710 0.300 ;
        RECT  1.300 -0.210 2.450 0.210 ;
        RECT  1.040 -0.210 1.300 0.310 ;
        RECT  0.260 -0.210 1.040 0.210 ;
        RECT  0.090 -0.210 0.260 0.520 ;
        RECT  0.000 -0.210 0.090 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.095 2.310 7.560 2.730 ;
        RECT  6.925 2.195 7.095 2.730 ;
        RECT  6.615 2.310 6.925 2.730 ;
        RECT  6.445 2.115 6.615 2.730 ;
        RECT  5.785 2.310 6.445 2.730 ;
        RECT  5.615 2.080 5.785 2.730 ;
        RECT  4.740 2.310 5.615 2.730 ;
        RECT  4.570 1.995 4.740 2.730 ;
        RECT  4.060 2.310 4.570 2.730 ;
        RECT  3.800 2.220 4.060 2.730 ;
        RECT  2.770 2.310 3.800 2.730 ;
        RECT  2.650 1.975 2.770 2.730 ;
        RECT  1.300 2.310 2.650 2.730 ;
        RECT  1.040 2.040 1.300 2.730 ;
        RECT  0.265 2.310 1.040 2.730 ;
        RECT  0.095 1.925 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  7.025 1.000 7.230 1.260 ;
        RECT  6.905 0.400 7.025 1.860 ;
        RECT  6.330 0.400 6.905 0.520 ;
        RECT  6.225 1.740 6.905 1.860 ;
        RECT  6.230 0.860 6.350 1.520 ;
        RECT  5.220 0.860 6.230 0.980 ;
        RECT  6.055 1.740 6.225 1.910 ;
        RECT  5.690 1.740 6.055 1.860 ;
        RECT  5.720 0.620 5.860 0.740 ;
        RECT  5.600 0.380 5.720 0.740 ;
        RECT  5.570 1.280 5.690 1.860 ;
        RECT  4.345 0.380 5.600 0.500 ;
        RECT  4.980 1.985 5.440 2.105 ;
        RECT  5.100 0.620 5.220 1.865 ;
        RECT  4.900 0.620 5.100 0.740 ;
        RECT  4.860 0.860 4.980 2.105 ;
        RECT  3.250 1.720 4.860 1.840 ;
        RECT  4.730 0.620 4.775 0.740 ;
        RECT  4.605 0.620 4.730 1.600 ;
        RECT  4.515 0.620 4.605 0.790 ;
        RECT  4.365 1.480 4.605 1.600 ;
        RECT  3.925 0.670 4.515 0.790 ;
        RECT  4.365 1.100 4.485 1.360 ;
        RECT  4.170 1.210 4.365 1.360 ;
        RECT  4.175 0.380 4.345 0.550 ;
        RECT  3.010 1.960 4.220 2.080 ;
        RECT  4.050 1.210 4.170 1.600 ;
        RECT  3.670 1.480 4.050 1.600 ;
        RECT  3.805 0.490 3.925 0.790 ;
        RECT  3.430 0.490 3.805 0.610 ;
        RECT  3.550 0.730 3.670 1.600 ;
        RECT  2.865 1.165 3.550 1.285 ;
        RECT  3.410 1.480 3.550 1.600 ;
        RECT  3.310 0.490 3.430 1.045 ;
        RECT  2.715 0.925 3.310 1.045 ;
        RECT  3.130 1.405 3.250 1.840 ;
        RECT  3.020 0.635 3.190 0.805 ;
        RECT  2.475 1.405 3.130 1.525 ;
        RECT  2.945 0.350 3.115 0.470 ;
        RECT  2.475 0.685 3.020 0.805 ;
        RECT  2.890 1.645 3.010 2.080 ;
        RECT  2.825 0.350 2.945 0.540 ;
        RECT  2.340 1.645 2.890 1.765 ;
        RECT  2.095 0.420 2.825 0.540 ;
        RECT  2.595 0.925 2.715 1.285 ;
        RECT  2.355 0.685 2.475 1.525 ;
        RECT  2.275 1.025 2.355 1.285 ;
        RECT  2.150 1.645 2.340 2.050 ;
        RECT  2.150 0.660 2.235 0.830 ;
        RECT  2.080 0.660 2.150 2.050 ;
        RECT  1.925 0.335 2.095 0.540 ;
        RECT  2.030 0.660 2.080 1.765 ;
        RECT  1.790 0.670 1.910 2.040 ;
        RECT  1.755 0.670 1.790 0.790 ;
        RECT  1.715 1.800 1.790 2.040 ;
        RECT  1.635 0.430 1.755 0.790 ;
        RECT  0.600 1.800 1.715 1.920 ;
        RECT  1.550 0.950 1.670 1.470 ;
        RECT  0.670 0.430 1.635 0.550 ;
        RECT  1.400 0.950 1.550 1.070 ;
        RECT  1.280 0.690 1.400 1.070 ;
        RECT  0.555 0.690 1.280 0.810 ;
        RECT  0.410 0.390 0.670 0.550 ;
        RECT  0.480 1.800 0.600 2.060 ;
        RECT  0.505 0.690 0.555 0.950 ;
        RECT  0.505 1.495 0.555 1.665 ;
        RECT  0.385 0.690 0.505 1.665 ;
    END
END SDFFSX1AD
MACRO SDFFSX2AD
    CLASS CORE ;
    FOREIGN SDFFSX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.910 1.100 6.090 1.620 ;
        RECT  5.840 1.360 5.910 1.620 ;
        END
        AntennaGateArea 0.101 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.965 1.580 1.430 1.700 ;
        RECT  0.965 0.930 1.130 1.070 ;
        RECT  0.845 0.930 0.965 1.700 ;
        RECT  0.630 1.145 0.845 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.265 1.280 ;
        RECT  0.070 1.020 0.210 1.655 ;
        END
        AntennaGateArea 0.103 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.770 0.735 6.930 1.545 ;
        RECT  6.585 0.735 6.770 0.905 ;
        RECT  6.585 1.375 6.770 1.545 ;
        END
        AntennaDiffArea 0.287 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.350 0.640 7.490 1.895 ;
        RECT  7.320 0.640 7.350 0.900 ;
        RECT  7.320 1.375 7.350 1.895 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.090 1.190 1.375 1.430 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.850 0.910 4.175 1.090 ;
        RECT  3.730 0.910 3.850 1.275 ;
        END
        AntennaGateArea 0.096 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.115 -0.210 7.560 0.210 ;
        RECT  6.945 -0.210 7.115 0.535 ;
        RECT  6.080 -0.210 6.945 0.210 ;
        RECT  5.820 -0.210 6.080 0.255 ;
        RECT  3.990 -0.210 5.820 0.210 ;
        RECT  3.730 -0.210 3.990 0.265 ;
        RECT  2.795 -0.210 3.730 0.210 ;
        RECT  2.535 -0.210 2.795 0.270 ;
        RECT  1.310 -0.210 2.535 0.210 ;
        RECT  1.050 -0.210 1.310 0.310 ;
        RECT  0.260 -0.210 1.050 0.210 ;
        RECT  0.090 -0.210 0.260 0.520 ;
        RECT  0.000 -0.210 0.090 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.115 2.310 7.560 2.730 ;
        RECT  6.945 1.980 7.115 2.730 ;
        RECT  6.485 2.310 6.945 2.730 ;
        RECT  6.315 2.225 6.485 2.730 ;
        RECT  5.745 2.310 6.315 2.730 ;
        RECT  5.575 2.080 5.745 2.730 ;
        RECT  4.670 2.310 5.575 2.730 ;
        RECT  4.500 2.020 4.670 2.730 ;
        RECT  4.010 2.310 4.500 2.730 ;
        RECT  3.750 2.220 4.010 2.730 ;
        RECT  2.730 2.310 3.750 2.730 ;
        RECT  2.610 2.005 2.730 2.730 ;
        RECT  1.300 2.310 2.610 2.730 ;
        RECT  1.040 2.060 1.300 2.730 ;
        RECT  0.255 2.310 1.040 2.730 ;
        RECT  0.085 1.900 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  7.200 1.000 7.230 1.260 ;
        RECT  7.080 1.000 7.200 1.860 ;
        RECT  6.455 1.740 7.080 1.860 ;
        RECT  6.335 0.330 6.455 1.860 ;
        RECT  6.165 1.740 6.335 1.860 ;
        RECT  6.070 0.375 6.190 0.980 ;
        RECT  5.995 1.740 6.165 1.910 ;
        RECT  5.160 0.860 6.070 0.980 ;
        RECT  5.650 1.740 5.995 1.860 ;
        RECT  5.560 0.620 5.700 0.740 ;
        RECT  5.530 1.295 5.650 1.860 ;
        RECT  5.440 0.380 5.560 0.740 ;
        RECT  4.285 0.380 5.440 0.500 ;
        RECT  4.910 1.985 5.410 2.105 ;
        RECT  5.040 0.620 5.160 1.735 ;
        RECT  4.820 0.620 5.040 0.740 ;
        RECT  4.790 0.860 4.910 2.105 ;
        RECT  4.780 0.860 4.790 1.830 ;
        RECT  3.210 1.710 4.780 1.830 ;
        RECT  4.660 0.620 4.690 0.740 ;
        RECT  4.540 0.620 4.660 1.590 ;
        RECT  4.430 0.620 4.540 0.790 ;
        RECT  4.335 1.470 4.540 1.590 ;
        RECT  3.865 0.670 4.430 0.790 ;
        RECT  4.300 1.090 4.420 1.350 ;
        RECT  4.110 1.230 4.300 1.350 ;
        RECT  4.115 0.380 4.285 0.550 ;
        RECT  2.970 1.960 4.190 2.080 ;
        RECT  3.990 1.230 4.110 1.590 ;
        RECT  3.610 1.470 3.990 1.590 ;
        RECT  3.745 0.385 3.865 0.790 ;
        RECT  3.370 0.385 3.745 0.505 ;
        RECT  3.490 0.625 3.610 1.590 ;
        RECT  2.900 1.175 3.490 1.295 ;
        RECT  3.370 1.470 3.490 1.590 ;
        RECT  3.250 0.385 3.370 1.055 ;
        RECT  2.720 0.935 3.250 1.055 ;
        RECT  3.090 1.520 3.210 1.830 ;
        RECT  2.960 0.645 3.130 0.815 ;
        RECT  2.415 1.520 3.090 1.640 ;
        RECT  2.005 0.390 3.055 0.510 ;
        RECT  2.850 1.760 2.970 2.080 ;
        RECT  2.415 0.695 2.960 0.815 ;
        RECT  2.265 1.760 2.850 1.880 ;
        RECT  2.600 0.935 2.720 1.400 ;
        RECT  2.295 0.695 2.415 1.640 ;
        RECT  2.225 1.025 2.295 1.285 ;
        RECT  2.145 1.760 2.265 1.945 ;
        RECT  2.100 0.645 2.175 0.815 ;
        RECT  2.100 1.435 2.145 1.945 ;
        RECT  2.095 0.645 2.100 1.945 ;
        RECT  2.025 0.645 2.095 1.880 ;
        RECT  1.980 0.645 2.025 1.555 ;
        RECT  1.835 0.335 2.005 0.510 ;
        RECT  1.740 0.670 1.860 2.085 ;
        RECT  1.700 0.670 1.740 0.790 ;
        RECT  0.625 1.820 1.740 1.940 ;
        RECT  1.580 0.430 1.700 0.790 ;
        RECT  1.500 0.920 1.620 1.440 ;
        RECT  0.670 0.430 1.580 0.550 ;
        RECT  1.400 0.920 1.500 1.040 ;
        RECT  1.280 0.690 1.400 1.040 ;
        RECT  0.555 0.690 1.280 0.810 ;
        RECT  0.410 0.390 0.670 0.550 ;
        RECT  0.455 1.820 0.625 2.015 ;
        RECT  0.505 0.690 0.555 0.950 ;
        RECT  0.505 1.470 0.555 1.640 ;
        RECT  0.385 0.690 0.505 1.640 ;
    END
END SDFFSX2AD
MACRO SDFFSX4AD
    CLASS CORE ;
    FOREIGN SDFFSX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.445 1.470 6.975 1.610 ;
        RECT  6.275 1.440 6.445 1.610 ;
        END
        AntennaGateArea 0.148 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.795 1.560 1.440 1.680 ;
        RECT  0.795 0.920 1.160 1.040 ;
        RECT  0.675 0.920 0.795 1.680 ;
        RECT  0.630 1.145 0.675 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.235 1.020 0.265 1.280 ;
        RECT  0.070 1.020 0.235 1.655 ;
        END
        AntennaGateArea 0.103 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.345 0.380 7.515 1.620 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.250 0.995 8.330 1.515 ;
        RECT  8.090 0.380 8.250 1.985 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.915 1.190 1.375 1.360 ;
        END
        AntennaGateArea 0.057 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.900 0.910 4.175 1.095 ;
        RECT  3.780 0.880 3.900 1.140 ;
        END
        AntennaGateArea 0.112 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.595 -0.210 8.680 0.210 ;
        RECT  8.425 -0.210 8.595 0.830 ;
        RECT  7.875 -0.210 8.425 0.210 ;
        RECT  7.705 -0.210 7.875 0.830 ;
        RECT  7.155 -0.210 7.705 0.210 ;
        RECT  6.985 -0.210 7.155 0.525 ;
        RECT  6.595 -0.210 6.985 0.210 ;
        RECT  6.425 -0.210 6.595 0.415 ;
        RECT  4.165 -0.210 6.425 0.210 ;
        RECT  3.905 -0.210 4.165 0.260 ;
        RECT  2.820 -0.210 3.905 0.210 ;
        RECT  2.560 -0.210 2.820 0.415 ;
        RECT  1.305 -0.210 2.560 0.210 ;
        RECT  1.045 -0.210 1.305 0.300 ;
        RECT  0.260 -0.210 1.045 0.210 ;
        RECT  0.120 -0.210 0.260 0.520 ;
        RECT  0.000 -0.210 0.120 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.595 2.310 8.680 2.730 ;
        RECT  8.425 1.650 8.595 2.730 ;
        RECT  7.875 2.310 8.425 2.730 ;
        RECT  7.705 1.985 7.875 2.730 ;
        RECT  7.155 2.310 7.705 2.730 ;
        RECT  6.985 1.985 7.155 2.730 ;
        RECT  6.335 2.310 6.985 2.730 ;
        RECT  6.165 2.065 6.335 2.730 ;
        RECT  5.095 2.310 6.165 2.730 ;
        RECT  4.925 2.065 5.095 2.730 ;
        RECT  4.690 2.310 4.925 2.730 ;
        RECT  4.520 2.065 4.690 2.730 ;
        RECT  4.050 2.310 4.520 2.730 ;
        RECT  3.790 1.950 4.050 2.730 ;
        RECT  2.750 2.310 3.790 2.730 ;
        RECT  2.630 2.025 2.750 2.730 ;
        RECT  1.255 2.310 2.630 2.730 ;
        RECT  1.085 2.050 1.255 2.730 ;
        RECT  0.240 2.310 1.085 2.730 ;
        RECT  0.120 1.880 0.240 2.730 ;
        RECT  0.000 2.310 0.120 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.680 2.520 ;
        LAYER M1 ;
        RECT  7.830 1.010 7.950 1.860 ;
        RECT  7.225 1.740 7.830 1.860 ;
        RECT  7.105 0.745 7.225 1.860 ;
        RECT  6.660 0.745 7.105 0.865 ;
        RECT  6.775 1.740 7.105 1.860 ;
        RECT  6.805 1.015 6.975 1.215 ;
        RECT  5.820 1.015 6.805 1.135 ;
        RECT  6.605 1.740 6.775 1.940 ;
        RECT  6.070 1.740 6.605 1.860 ;
        RECT  6.155 0.595 6.205 0.765 ;
        RECT  6.035 0.380 6.155 0.765 ;
        RECT  5.950 1.410 6.070 1.860 ;
        RECT  4.610 0.380 6.035 0.500 ;
        RECT  5.700 0.620 5.820 1.535 ;
        RECT  5.550 2.020 5.810 2.190 ;
        RECT  5.380 0.620 5.700 0.740 ;
        RECT  5.625 1.415 5.700 1.535 ;
        RECT  5.455 1.415 5.625 1.880 ;
        RECT  5.335 2.020 5.550 2.140 ;
        RECT  5.335 0.910 5.515 1.030 ;
        RECT  5.215 0.910 5.335 2.140 ;
        RECT  4.940 0.620 5.260 0.740 ;
        RECT  3.230 1.710 5.215 1.830 ;
        RECT  4.820 0.620 4.940 1.575 ;
        RECT  4.465 0.620 4.820 0.740 ;
        RECT  4.395 1.455 4.820 1.575 ;
        RECT  4.350 1.060 4.470 1.335 ;
        RECT  4.345 0.365 4.465 0.740 ;
        RECT  4.235 1.215 4.350 1.335 ;
        RECT  4.295 0.365 4.345 0.535 ;
        RECT  3.405 0.380 4.295 0.500 ;
        RECT  4.115 1.215 4.235 1.545 ;
        RECT  3.645 1.425 4.115 1.545 ;
        RECT  3.645 0.620 3.785 0.740 ;
        RECT  3.525 0.620 3.645 1.545 ;
        RECT  3.455 1.145 3.525 1.545 ;
        RECT  3.220 2.020 3.480 2.190 ;
        RECT  2.910 1.145 3.455 1.265 ;
        RECT  3.285 0.380 3.405 1.025 ;
        RECT  2.725 0.905 3.285 1.025 ;
        RECT  3.110 1.385 3.230 1.830 ;
        RECT  2.990 2.020 3.220 2.140 ;
        RECT  3.045 0.525 3.165 0.785 ;
        RECT  2.485 1.385 3.110 1.505 ;
        RECT  2.485 0.665 3.045 0.785 ;
        RECT  2.870 1.625 2.990 2.140 ;
        RECT  2.265 1.625 2.870 1.745 ;
        RECT  2.605 0.905 2.725 1.265 ;
        RECT  2.365 0.665 2.485 1.505 ;
        RECT  2.275 1.075 2.365 1.335 ;
        RECT  2.150 1.625 2.265 2.070 ;
        RECT  2.150 0.655 2.245 0.915 ;
        RECT  2.095 0.655 2.150 2.070 ;
        RECT  2.030 0.655 2.095 1.745 ;
        RECT  1.790 0.420 1.910 2.040 ;
        RECT  1.735 0.420 1.790 0.820 ;
        RECT  1.715 1.800 1.790 2.040 ;
        RECT  0.410 0.420 1.735 0.540 ;
        RECT  0.600 1.800 1.715 1.920 ;
        RECT  1.615 1.130 1.670 1.390 ;
        RECT  1.495 0.680 1.615 1.390 ;
        RECT  0.555 0.680 1.495 0.800 ;
        RECT  0.480 1.800 0.600 2.060 ;
        RECT  0.505 0.680 0.555 0.905 ;
        RECT  0.505 1.495 0.555 1.665 ;
        RECT  0.385 0.680 0.505 1.665 ;
    END
END SDFFSX4AD
MACRO SDFFSXLAD
    CLASS CORE ;
    FOREIGN SDFFSXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.910 1.100 6.090 1.620 ;
        END
        AntennaGateArea 0.081 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.995 1.560 1.430 1.680 ;
        RECT  0.995 0.930 1.160 1.070 ;
        RECT  0.875 0.930 0.995 1.680 ;
        RECT  0.630 1.145 0.875 1.375 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.020 0.265 1.280 ;
        RECT  0.070 1.020 0.210 1.655 ;
        END
        AntennaGateArea 0.103 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.670 0.690 6.780 0.950 ;
        RECT  6.670 1.330 6.780 1.590 ;
        RECT  6.510 0.690 6.670 1.590 ;
        END
        AntennaDiffArea 0.129 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.350 0.735 7.490 1.695 ;
        RECT  7.305 0.735 7.350 0.905 ;
        RECT  7.320 1.375 7.350 1.695 ;
        END
        AntennaDiffArea 0.143 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.115 1.190 1.415 1.430 ;
        END
        AntennaGateArea 0.055 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.925 0.910 4.175 1.090 ;
        RECT  3.805 0.910 3.925 1.275 ;
        END
        AntennaGateArea 0.089 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.265 -0.210 7.560 0.210 ;
        RECT  7.145 -0.210 7.265 0.420 ;
        RECT  6.240 -0.210 7.145 0.210 ;
        RECT  5.980 -0.210 6.240 0.310 ;
        RECT  4.005 -0.210 5.980 0.210 ;
        RECT  3.835 -0.210 4.005 0.370 ;
        RECT  2.710 -0.210 3.835 0.210 ;
        RECT  2.450 -0.210 2.710 0.300 ;
        RECT  1.300 -0.210 2.450 0.210 ;
        RECT  1.040 -0.210 1.300 0.310 ;
        RECT  0.260 -0.210 1.040 0.210 ;
        RECT  0.090 -0.210 0.260 0.520 ;
        RECT  0.000 -0.210 0.090 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.095 2.310 7.560 2.730 ;
        RECT  6.925 2.015 7.095 2.730 ;
        RECT  6.615 2.310 6.925 2.730 ;
        RECT  6.445 1.980 6.615 2.730 ;
        RECT  5.785 2.310 6.445 2.730 ;
        RECT  5.615 2.080 5.785 2.730 ;
        RECT  4.740 2.310 5.615 2.730 ;
        RECT  4.570 1.995 4.740 2.730 ;
        RECT  4.060 2.310 4.570 2.730 ;
        RECT  3.800 2.220 4.060 2.730 ;
        RECT  2.770 2.310 3.800 2.730 ;
        RECT  2.650 1.975 2.770 2.730 ;
        RECT  1.300 2.310 2.650 2.730 ;
        RECT  1.040 2.040 1.300 2.730 ;
        RECT  0.265 2.310 1.040 2.730 ;
        RECT  0.095 1.925 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  7.025 1.000 7.230 1.260 ;
        RECT  6.905 0.400 7.025 1.860 ;
        RECT  6.330 0.400 6.905 0.520 ;
        RECT  6.225 1.740 6.905 1.860 ;
        RECT  6.230 0.860 6.350 1.520 ;
        RECT  5.220 0.860 6.230 0.980 ;
        RECT  6.055 1.740 6.225 1.910 ;
        RECT  5.690 1.740 6.055 1.860 ;
        RECT  5.720 0.620 5.860 0.740 ;
        RECT  5.600 0.380 5.720 0.740 ;
        RECT  5.570 1.280 5.690 1.860 ;
        RECT  4.345 0.380 5.600 0.500 ;
        RECT  4.980 1.985 5.440 2.105 ;
        RECT  5.100 0.620 5.220 1.865 ;
        RECT  4.900 0.620 5.100 0.740 ;
        RECT  4.860 0.860 4.980 2.105 ;
        RECT  3.250 1.720 4.860 1.840 ;
        RECT  4.730 0.620 4.775 0.740 ;
        RECT  4.605 0.620 4.730 1.600 ;
        RECT  4.515 0.620 4.605 0.790 ;
        RECT  4.365 1.480 4.605 1.600 ;
        RECT  3.925 0.670 4.515 0.790 ;
        RECT  4.365 1.100 4.485 1.360 ;
        RECT  4.170 1.210 4.365 1.360 ;
        RECT  4.175 0.380 4.345 0.550 ;
        RECT  3.010 1.960 4.220 2.080 ;
        RECT  4.050 1.210 4.170 1.600 ;
        RECT  3.670 1.480 4.050 1.600 ;
        RECT  3.805 0.490 3.925 0.790 ;
        RECT  3.430 0.490 3.805 0.610 ;
        RECT  3.550 0.730 3.670 1.600 ;
        RECT  2.865 1.165 3.550 1.285 ;
        RECT  3.410 1.480 3.550 1.600 ;
        RECT  3.310 0.490 3.430 1.045 ;
        RECT  2.715 0.925 3.310 1.045 ;
        RECT  3.130 1.405 3.250 1.840 ;
        RECT  3.020 0.635 3.190 0.805 ;
        RECT  2.475 1.405 3.130 1.525 ;
        RECT  2.945 0.350 3.115 0.470 ;
        RECT  2.475 0.685 3.020 0.805 ;
        RECT  2.890 1.645 3.010 2.080 ;
        RECT  2.825 0.350 2.945 0.540 ;
        RECT  2.340 1.645 2.890 1.765 ;
        RECT  2.095 0.420 2.825 0.540 ;
        RECT  2.595 0.925 2.715 1.285 ;
        RECT  2.355 0.685 2.475 1.525 ;
        RECT  2.275 1.025 2.355 1.285 ;
        RECT  2.150 1.645 2.340 2.050 ;
        RECT  2.150 0.660 2.235 0.830 ;
        RECT  2.080 0.660 2.150 2.050 ;
        RECT  1.925 0.335 2.095 0.540 ;
        RECT  2.030 0.660 2.080 1.765 ;
        RECT  1.790 0.670 1.910 2.040 ;
        RECT  1.755 0.670 1.790 0.790 ;
        RECT  1.715 1.800 1.790 2.040 ;
        RECT  1.635 0.430 1.755 0.790 ;
        RECT  0.600 1.800 1.715 1.920 ;
        RECT  1.550 0.950 1.670 1.470 ;
        RECT  0.670 0.430 1.635 0.550 ;
        RECT  1.400 0.950 1.550 1.070 ;
        RECT  1.280 0.690 1.400 1.070 ;
        RECT  0.555 0.690 1.280 0.810 ;
        RECT  0.410 0.390 0.670 0.550 ;
        RECT  0.480 1.800 0.600 2.060 ;
        RECT  0.505 0.690 0.555 0.950 ;
        RECT  0.505 1.495 0.555 1.665 ;
        RECT  0.385 0.690 0.505 1.665 ;
    END
END SDFFSXLAD
MACRO SDFFTRX1AD
    CLASS CORE ;
    FOREIGN SDFFTRX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 0.890 2.215 1.060 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.970 2.460 2.090 ;
        RECT  1.185 1.970 1.440 2.190 ;
        RECT  1.065 1.730 1.185 2.190 ;
        RECT  0.610 1.730 1.065 1.890 ;
        RECT  0.350 1.330 0.610 1.890 ;
        END
        AntennaGateArea 0.134 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.510 2.495 1.125 ;
        RECT  2.265 0.510 2.345 0.770 ;
        RECT  1.920 0.510 2.265 0.630 ;
        RECT  1.800 0.380 1.920 0.630 ;
        RECT  1.055 0.380 1.800 0.500 ;
        RECT  0.935 0.380 1.055 0.830 ;
        RECT  0.780 0.710 0.935 0.830 ;
        RECT  0.660 0.710 0.780 0.970 ;
        END
        AntennaGateArea 0.055 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.145 0.705 7.330 1.530 ;
        RECT  7.060 1.145 7.145 1.530 ;
        END
        AntennaDiffArea 0.181 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.010 0.645 8.050 1.530 ;
        RECT  7.890 0.645 8.010 1.860 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 1.330 1.145 1.610 ;
        END
        AntennaGateArea 0.065 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.905 1.110 3.335 1.330 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.675 -0.210 8.120 0.210 ;
        RECT  7.505 -0.210 7.675 0.825 ;
        RECT  6.580 -0.210 7.505 0.210 ;
        RECT  6.320 -0.210 6.580 0.730 ;
        RECT  5.155 -0.210 6.320 0.210 ;
        RECT  4.895 -0.210 5.155 0.300 ;
        RECT  3.285 -0.210 4.895 0.210 ;
        RECT  3.025 -0.210 3.285 0.635 ;
        RECT  2.210 -0.210 3.025 0.210 ;
        RECT  2.040 -0.210 2.210 0.390 ;
        RECT  0.655 -0.210 2.040 0.210 ;
        RECT  0.485 -0.210 0.655 0.590 ;
        RECT  0.000 -0.210 0.485 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.655 2.310 8.120 2.730 ;
        RECT  7.485 1.905 7.655 2.730 ;
        RECT  6.695 2.310 7.485 2.730 ;
        RECT  6.525 2.220 6.695 2.730 ;
        RECT  5.095 2.310 6.525 2.730 ;
        RECT  4.925 1.785 5.095 2.730 ;
        RECT  3.500 2.310 4.925 2.730 ;
        RECT  3.240 2.200 3.500 2.730 ;
        RECT  2.270 2.310 3.240 2.730 ;
        RECT  2.010 2.230 2.270 2.730 ;
        RECT  0.885 2.310 2.010 2.730 ;
        RECT  0.455 2.095 0.885 2.730 ;
        RECT  0.000 2.310 0.455 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.120 2.520 ;
        LAYER M1 ;
        RECT  7.650 1.010 7.770 1.780 ;
        RECT  6.990 1.650 7.650 1.780 ;
        RECT  6.905 1.650 6.990 2.100 ;
        RECT  6.785 0.540 6.905 2.100 ;
        RECT  6.405 1.980 6.785 2.100 ;
        RECT  6.545 1.025 6.665 1.545 ;
        RECT  6.420 0.850 6.545 1.850 ;
        RECT  5.890 0.850 6.420 0.970 ;
        RECT  5.600 1.730 6.420 1.850 ;
        RECT  6.235 1.980 6.405 2.185 ;
        RECT  5.820 1.175 6.080 1.570 ;
        RECT  5.770 0.540 5.890 0.970 ;
        RECT  5.650 1.175 5.820 1.300 ;
        RECT  5.530 0.420 5.650 1.300 ;
        RECT  4.730 0.420 5.530 0.540 ;
        RECT  5.410 1.450 5.480 1.970 ;
        RECT  5.290 0.660 5.410 1.970 ;
        RECT  5.260 0.660 5.290 0.920 ;
        RECT  4.900 0.800 5.260 0.920 ;
        RECT  5.050 1.040 5.170 1.515 ;
        RECT  4.510 1.395 5.050 1.515 ;
        RECT  4.780 0.800 4.900 1.265 ;
        RECT  4.640 1.145 4.780 1.265 ;
        RECT  4.610 0.380 4.730 0.540 ;
        RECT  3.830 0.380 4.610 0.500 ;
        RECT  4.390 0.640 4.510 2.125 ;
        RECT  4.310 0.640 4.390 0.810 ;
        RECT  4.295 1.925 4.390 2.125 ;
        RECT  4.045 0.640 4.165 2.095 ;
        RECT  3.950 0.640 4.045 0.810 ;
        RECT  3.935 1.740 4.045 2.095 ;
        RECT  2.940 1.740 3.935 1.860 ;
        RECT  3.830 1.070 3.925 1.555 ;
        RECT  3.710 0.380 3.830 1.555 ;
        RECT  3.430 0.490 3.710 0.660 ;
        RECT  3.675 1.385 3.710 1.555 ;
        RECT  3.470 0.780 3.590 1.300 ;
        RECT  2.850 0.780 3.470 0.900 ;
        RECT  2.780 1.450 3.210 1.570 ;
        RECT  2.680 1.710 2.940 1.910 ;
        RECT  2.780 0.490 2.850 0.900 ;
        RECT  2.660 0.490 2.780 1.570 ;
        RECT  2.040 1.710 2.680 1.830 ;
        RECT  1.920 1.180 2.040 1.830 ;
        RECT  1.680 1.180 1.920 1.300 ;
        RECT  1.355 1.710 1.920 1.830 ;
        RECT  1.440 1.420 1.770 1.540 ;
        RECT  1.560 0.620 1.680 1.300 ;
        RECT  1.330 0.620 1.560 0.740 ;
        RECT  1.315 0.880 1.440 1.540 ;
        RECT  1.180 0.880 1.315 1.210 ;
        RECT  0.230 1.090 1.180 1.210 ;
        RECT  0.110 0.400 0.230 1.810 ;
    END
END SDFFTRX1AD
MACRO SDFFTRX2AD
    CLASS CORE ;
    FOREIGN SDFFTRX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 0.890 2.215 1.060 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.970 2.460 2.090 ;
        RECT  1.185 1.970 1.440 2.190 ;
        RECT  1.065 1.730 1.185 2.190 ;
        RECT  0.610 1.730 1.065 1.890 ;
        RECT  0.350 1.330 0.610 1.890 ;
        END
        AntennaGateArea 0.133 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.510 2.495 1.125 ;
        RECT  2.265 0.510 2.345 0.770 ;
        RECT  1.920 0.510 2.265 0.630 ;
        RECT  1.800 0.380 1.920 0.630 ;
        RECT  1.055 0.380 1.800 0.500 ;
        RECT  0.935 0.380 1.055 0.830 ;
        RECT  0.780 0.710 0.935 0.830 ;
        RECT  0.660 0.710 0.780 0.970 ;
        END
        AntennaGateArea 0.055 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.320 0.760 7.360 0.880 ;
        RECT  7.070 0.760 7.320 1.555 ;
        END
        AntennaDiffArea 0.322 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.010 0.645 8.050 1.530 ;
        RECT  7.890 0.395 8.010 1.950 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 1.330 1.145 1.610 ;
        END
        AntennaGateArea 0.064 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.905 1.110 3.335 1.330 ;
        END
        AntennaGateArea 0.077 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.720 -0.210 8.120 0.210 ;
        RECT  7.460 -0.210 7.720 0.390 ;
        RECT  6.725 -0.210 7.460 0.210 ;
        RECT  6.715 -0.210 6.725 0.220 ;
        RECT  6.455 -0.210 6.715 0.240 ;
        RECT  5.180 -0.210 6.455 0.210 ;
        RECT  4.920 -0.210 5.180 0.260 ;
        RECT  3.285 -0.210 4.920 0.210 ;
        RECT  3.025 -0.210 3.285 0.635 ;
        RECT  2.210 -0.210 3.025 0.210 ;
        RECT  2.040 -0.210 2.210 0.390 ;
        RECT  0.655 -0.210 2.040 0.210 ;
        RECT  0.485 -0.210 0.655 0.590 ;
        RECT  0.000 -0.210 0.485 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.655 2.310 8.120 2.730 ;
        RECT  7.485 1.975 7.655 2.730 ;
        RECT  6.655 2.310 7.485 2.730 ;
        RECT  6.485 2.220 6.655 2.730 ;
        RECT  5.180 2.310 6.485 2.730 ;
        RECT  4.920 2.210 5.180 2.730 ;
        RECT  3.500 2.310 4.920 2.730 ;
        RECT  3.240 2.200 3.500 2.730 ;
        RECT  2.270 2.310 3.240 2.730 ;
        RECT  2.010 2.230 2.270 2.730 ;
        RECT  0.885 2.310 2.010 2.730 ;
        RECT  0.455 2.095 0.885 2.730 ;
        RECT  0.000 2.310 0.455 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.120 2.520 ;
        LAYER M1 ;
        RECT  7.650 0.520 7.770 1.800 ;
        RECT  6.950 0.520 7.650 0.640 ;
        RECT  6.980 1.680 7.650 1.800 ;
        RECT  6.965 1.680 6.980 1.945 ;
        RECT  6.845 1.680 6.965 1.950 ;
        RECT  6.830 0.480 6.950 0.740 ;
        RECT  6.370 1.830 6.845 1.950 ;
        RECT  6.680 0.885 6.800 1.405 ;
        RECT  6.350 1.095 6.680 1.215 ;
        RECT  6.250 1.830 6.370 2.090 ;
        RECT  6.230 0.910 6.350 1.710 ;
        RECT  5.995 0.910 6.230 1.030 ;
        RECT  5.730 1.590 6.230 1.710 ;
        RECT  5.755 1.310 6.110 1.430 ;
        RECT  5.760 2.070 6.110 2.190 ;
        RECT  5.875 0.420 5.995 1.030 ;
        RECT  5.640 1.970 5.760 2.190 ;
        RECT  5.635 0.380 5.755 1.430 ;
        RECT  4.700 1.970 5.640 2.090 ;
        RECT  3.830 0.380 5.635 0.500 ;
        RECT  5.490 0.620 5.515 0.790 ;
        RECT  5.370 0.620 5.490 1.710 ;
        RECT  5.345 0.620 5.370 0.790 ;
        RECT  4.870 0.670 5.345 0.790 ;
        RECT  5.130 1.040 5.250 1.620 ;
        RECT  4.440 1.500 5.130 1.620 ;
        RECT  4.750 0.670 4.870 1.315 ;
        RECT  4.580 1.890 4.700 2.150 ;
        RECT  4.440 0.635 4.480 0.805 ;
        RECT  4.320 0.635 4.440 2.140 ;
        RECT  4.310 0.635 4.320 0.805 ;
        RECT  4.045 0.635 4.165 2.095 ;
        RECT  3.950 0.635 4.045 0.805 ;
        RECT  3.935 1.740 4.045 2.095 ;
        RECT  2.940 1.740 3.935 1.860 ;
        RECT  3.830 1.070 3.925 1.555 ;
        RECT  3.710 0.380 3.830 1.555 ;
        RECT  3.430 0.490 3.710 0.660 ;
        RECT  3.675 1.385 3.710 1.555 ;
        RECT  3.470 0.780 3.590 1.300 ;
        RECT  2.850 0.780 3.470 0.900 ;
        RECT  2.780 1.450 3.210 1.570 ;
        RECT  2.680 1.710 2.940 1.910 ;
        RECT  2.780 0.490 2.850 0.900 ;
        RECT  2.660 0.490 2.780 1.570 ;
        RECT  2.040 1.710 2.680 1.830 ;
        RECT  1.920 1.180 2.040 1.830 ;
        RECT  1.680 1.180 1.920 1.300 ;
        RECT  1.355 1.710 1.920 1.830 ;
        RECT  1.440 1.420 1.770 1.540 ;
        RECT  1.560 0.620 1.680 1.300 ;
        RECT  1.330 0.620 1.560 0.740 ;
        RECT  1.315 0.880 1.440 1.540 ;
        RECT  1.180 0.880 1.315 1.210 ;
        RECT  0.230 1.090 1.180 1.210 ;
        RECT  0.110 0.400 0.230 1.810 ;
    END
END SDFFTRX2AD
MACRO SDFFTRX4AD
    CLASS CORE ;
    FOREIGN SDFFTRX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 0.890 2.215 1.060 ;
        END
        AntennaGateArea 0.055 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.445 1.970 2.460 2.090 ;
        RECT  1.305 1.970 1.445 2.190 ;
        RECT  1.185 1.730 1.305 2.190 ;
        RECT  0.610 1.730 1.185 1.890 ;
        RECT  0.350 1.330 0.610 1.890 ;
        END
        AntennaGateArea 0.162 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.510 2.495 1.125 ;
        RECT  2.265 0.510 2.345 0.770 ;
        RECT  1.920 0.510 2.265 0.630 ;
        RECT  1.800 0.380 1.920 0.630 ;
        RECT  1.055 0.380 1.800 0.500 ;
        RECT  0.935 0.380 1.055 0.970 ;
        RECT  0.560 0.850 0.935 0.970 ;
        END
        AntennaGateArea 0.078 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.745 0.450 8.960 1.530 ;
        RECT  8.700 1.145 8.745 1.530 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.590 0.405 9.730 1.945 ;
        RECT  9.465 0.405 9.590 0.835 ;
        RECT  9.490 1.425 9.590 1.945 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.815 2.070 1.065 2.190 ;
        RECT  0.585 2.030 0.815 2.190 ;
        END
        AntennaGateArea 0.105 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.905 1.110 3.335 1.330 ;
        END
        AntennaGateArea 0.113 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.970 -0.210 10.080 0.210 ;
        RECT  9.850 -0.210 9.970 0.815 ;
        RECT  9.275 -0.210 9.850 0.210 ;
        RECT  9.105 -0.210 9.275 0.770 ;
        RECT  8.530 -0.210 9.105 0.210 ;
        RECT  8.270 -0.210 8.530 0.260 ;
        RECT  7.880 -0.210 8.270 0.210 ;
        RECT  7.620 -0.210 7.880 0.450 ;
        RECT  6.000 -0.210 7.620 0.210 ;
        RECT  5.740 -0.210 6.000 0.260 ;
        RECT  5.235 -0.210 5.740 0.210 ;
        RECT  4.975 -0.210 5.235 0.260 ;
        RECT  3.285 -0.210 4.975 0.210 ;
        RECT  3.025 -0.210 3.285 0.635 ;
        RECT  2.210 -0.210 3.025 0.210 ;
        RECT  2.040 -0.210 2.210 0.390 ;
        RECT  0.655 -0.210 2.040 0.210 ;
        RECT  0.485 -0.210 0.655 0.715 ;
        RECT  0.000 -0.210 0.485 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.970 2.310 10.080 2.730 ;
        RECT  9.850 1.735 9.970 2.730 ;
        RECT  9.275 2.310 9.850 2.730 ;
        RECT  9.105 1.975 9.275 2.730 ;
        RECT  8.485 2.310 9.105 2.730 ;
        RECT  8.315 2.175 8.485 2.730 ;
        RECT  7.905 2.310 8.315 2.730 ;
        RECT  7.735 2.175 7.905 2.730 ;
        RECT  6.000 2.310 7.735 2.730 ;
        RECT  5.740 2.240 6.000 2.730 ;
        RECT  5.240 2.310 5.740 2.730 ;
        RECT  4.980 2.240 5.240 2.730 ;
        RECT  3.590 2.310 4.980 2.730 ;
        RECT  3.330 2.200 3.590 2.730 ;
        RECT  2.270 2.310 3.330 2.730 ;
        RECT  2.010 2.230 2.270 2.730 ;
        RECT  0.465 2.310 2.010 2.730 ;
        RECT  0.295 2.095 0.465 2.730 ;
        RECT  0.000 2.310 0.295 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.080 2.520 ;
        LAYER M1 ;
        RECT  9.360 1.010 9.460 1.270 ;
        RECT  9.240 1.010 9.360 1.780 ;
        RECT  8.285 1.650 9.240 1.780 ;
        RECT  8.160 0.640 8.285 2.020 ;
        RECT  8.070 0.640 8.160 0.900 ;
        RECT  8.115 1.730 8.160 2.020 ;
        RECT  7.485 1.900 8.115 2.020 ;
        RECT  7.935 1.155 8.040 1.415 ;
        RECT  7.815 0.850 7.935 1.740 ;
        RECT  7.195 0.850 7.815 0.970 ;
        RECT  7.125 1.620 7.815 1.740 ;
        RECT  7.175 1.175 7.435 1.460 ;
        RECT  7.075 0.650 7.195 0.970 ;
        RECT  6.955 1.175 7.175 1.300 ;
        RECT  7.005 1.620 7.125 1.880 ;
        RECT  6.265 1.760 7.005 1.880 ;
        RECT  6.835 0.380 6.955 1.300 ;
        RECT  6.010 1.520 6.885 1.640 ;
        RECT  3.830 0.380 6.835 0.500 ;
        RECT  6.195 0.920 6.835 1.180 ;
        RECT  6.010 0.650 6.645 0.770 ;
        RECT  6.120 2.000 6.290 2.190 ;
        RECT  4.700 2.000 6.120 2.120 ;
        RECT  5.890 0.650 6.010 1.640 ;
        RECT  4.875 0.650 5.890 0.770 ;
        RECT  5.620 1.395 5.890 1.515 ;
        RECT  5.240 1.085 5.695 1.255 ;
        RECT  5.360 1.395 5.620 1.800 ;
        RECT  5.120 1.085 5.240 1.620 ;
        RECT  4.440 1.500 5.120 1.620 ;
        RECT  4.755 0.650 4.875 1.335 ;
        RECT  4.580 1.895 4.700 2.155 ;
        RECT  4.440 0.635 4.480 0.805 ;
        RECT  4.320 0.635 4.440 2.140 ;
        RECT  4.310 0.635 4.320 0.805 ;
        RECT  4.045 0.635 4.165 2.095 ;
        RECT  3.960 0.635 4.045 0.895 ;
        RECT  3.935 1.725 4.045 2.095 ;
        RECT  2.940 1.725 3.935 1.845 ;
        RECT  3.830 1.070 3.925 1.555 ;
        RECT  3.710 0.380 3.830 1.555 ;
        RECT  3.430 0.490 3.710 0.660 ;
        RECT  3.675 1.385 3.710 1.555 ;
        RECT  3.470 0.780 3.590 1.300 ;
        RECT  2.880 0.780 3.470 0.900 ;
        RECT  2.780 1.450 3.210 1.570 ;
        RECT  2.680 1.725 2.940 1.910 ;
        RECT  2.780 0.490 2.880 0.900 ;
        RECT  2.660 0.490 2.780 1.570 ;
        RECT  2.040 1.725 2.680 1.845 ;
        RECT  1.920 1.180 2.040 1.845 ;
        RECT  1.680 1.180 1.920 1.300 ;
        RECT  1.595 1.725 1.920 1.845 ;
        RECT  1.440 1.420 1.760 1.540 ;
        RECT  1.560 0.620 1.680 1.300 ;
        RECT  1.425 1.675 1.595 1.845 ;
        RECT  1.330 0.620 1.560 0.740 ;
        RECT  1.315 0.880 1.440 1.540 ;
        RECT  1.180 0.880 1.315 1.210 ;
        RECT  0.230 1.090 1.180 1.210 ;
        RECT  0.110 0.500 0.230 1.810 ;
    END
END SDFFTRX4AD
MACRO SDFFTRXLAD
    CLASS CORE ;
    FOREIGN SDFFTRXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 0.890 2.215 1.060 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.970 2.460 2.090 ;
        RECT  1.185 1.970 1.440 2.190 ;
        RECT  1.065 1.730 1.185 2.190 ;
        RECT  0.610 1.730 1.065 1.890 ;
        RECT  0.350 1.330 0.610 1.890 ;
        END
        AntennaGateArea 0.134 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.345 0.510 2.495 1.125 ;
        RECT  2.265 0.510 2.345 0.770 ;
        RECT  1.920 0.510 2.265 0.630 ;
        RECT  1.800 0.380 1.920 0.630 ;
        RECT  1.055 0.380 1.800 0.500 ;
        RECT  0.935 0.380 1.055 0.830 ;
        RECT  0.780 0.710 0.935 0.830 ;
        RECT  0.660 0.710 0.780 0.970 ;
        END
        AntennaGateArea 0.055 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.180 1.145 7.210 1.375 ;
        RECT  7.060 0.830 7.180 1.375 ;
        RECT  6.940 0.690 7.060 0.950 ;
        RECT  6.940 1.145 7.060 1.590 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.650 0.715 7.770 1.685 ;
        RECT  7.585 0.715 7.650 0.885 ;
        RECT  7.610 1.425 7.650 1.685 ;
        END
        AntennaDiffArea 0.143 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 1.330 1.145 1.610 ;
        END
        AntennaGateArea 0.065 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.905 1.110 3.335 1.330 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.375 -0.210 7.840 0.210 ;
        RECT  7.205 -0.210 7.375 0.475 ;
        RECT  6.580 -0.210 7.205 0.210 ;
        RECT  6.320 -0.210 6.580 0.540 ;
        RECT  5.125 -0.210 6.320 0.210 ;
        RECT  4.865 -0.210 5.125 0.300 ;
        RECT  3.285 -0.210 4.865 0.210 ;
        RECT  3.025 -0.210 3.285 0.635 ;
        RECT  2.210 -0.210 3.025 0.210 ;
        RECT  2.040 -0.210 2.210 0.390 ;
        RECT  0.655 -0.210 2.040 0.210 ;
        RECT  0.485 -0.210 0.655 0.590 ;
        RECT  0.000 -0.210 0.485 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.465 2.310 7.840 2.730 ;
        RECT  7.295 2.005 7.465 2.730 ;
        RECT  6.655 2.310 7.295 2.730 ;
        RECT  6.395 2.270 6.655 2.730 ;
        RECT  5.095 2.310 6.395 2.730 ;
        RECT  4.925 1.785 5.095 2.730 ;
        RECT  3.500 2.310 4.925 2.730 ;
        RECT  3.240 2.200 3.500 2.730 ;
        RECT  2.270 2.310 3.240 2.730 ;
        RECT  2.010 2.230 2.270 2.730 ;
        RECT  0.885 2.310 2.010 2.730 ;
        RECT  0.455 2.095 0.885 2.730 ;
        RECT  0.000 2.310 0.455 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.840 2.520 ;
        LAYER M1 ;
        RECT  7.490 1.010 7.520 1.270 ;
        RECT  7.370 1.010 7.490 1.885 ;
        RECT  6.990 1.755 7.370 1.885 ;
        RECT  6.820 1.755 6.990 2.130 ;
        RECT  6.820 0.420 6.975 0.540 ;
        RECT  6.700 0.420 6.820 2.130 ;
        RECT  6.180 2.010 6.700 2.130 ;
        RECT  6.545 1.020 6.580 1.280 ;
        RECT  6.420 0.850 6.545 1.850 ;
        RECT  5.880 0.850 6.420 0.970 ;
        RECT  5.600 1.730 6.420 1.850 ;
        RECT  5.810 1.175 6.070 1.570 ;
        RECT  5.760 0.350 5.880 0.970 ;
        RECT  5.640 1.175 5.810 1.300 ;
        RECT  5.520 0.420 5.640 1.300 ;
        RECT  4.730 0.420 5.520 0.540 ;
        RECT  5.400 1.635 5.455 1.805 ;
        RECT  5.280 0.660 5.400 1.805 ;
        RECT  5.250 0.660 5.280 0.920 ;
        RECT  4.900 0.800 5.250 0.920 ;
        RECT  5.040 1.040 5.160 1.515 ;
        RECT  4.510 1.395 5.040 1.515 ;
        RECT  4.780 0.800 4.900 1.265 ;
        RECT  4.640 1.145 4.780 1.265 ;
        RECT  4.610 0.380 4.730 0.540 ;
        RECT  3.830 0.380 4.610 0.500 ;
        RECT  4.390 0.640 4.510 2.050 ;
        RECT  4.310 0.640 4.390 0.810 ;
        RECT  4.295 1.880 4.390 2.050 ;
        RECT  4.045 0.640 4.165 2.095 ;
        RECT  3.950 0.640 4.045 0.810 ;
        RECT  3.935 1.740 4.045 2.095 ;
        RECT  2.940 1.740 3.935 1.860 ;
        RECT  3.830 1.070 3.925 1.555 ;
        RECT  3.710 0.380 3.830 1.555 ;
        RECT  3.430 0.490 3.710 0.660 ;
        RECT  3.675 1.385 3.710 1.555 ;
        RECT  3.470 0.780 3.590 1.300 ;
        RECT  2.850 0.780 3.470 0.900 ;
        RECT  2.780 1.450 3.210 1.570 ;
        RECT  2.680 1.710 2.940 1.910 ;
        RECT  2.780 0.490 2.850 0.900 ;
        RECT  2.660 0.490 2.780 1.570 ;
        RECT  2.040 1.710 2.680 1.830 ;
        RECT  1.920 1.180 2.040 1.830 ;
        RECT  1.680 1.180 1.920 1.300 ;
        RECT  1.355 1.710 1.920 1.830 ;
        RECT  1.440 1.420 1.770 1.540 ;
        RECT  1.560 0.620 1.680 1.300 ;
        RECT  1.330 0.620 1.560 0.740 ;
        RECT  1.315 0.880 1.440 1.540 ;
        RECT  1.180 0.880 1.315 1.210 ;
        RECT  0.230 1.090 1.180 1.210 ;
        RECT  0.110 0.400 0.230 1.810 ;
    END
END SDFFTRXLAD
MACRO SDFFX1AD
    CLASS CORE ;
    FOREIGN SDFFX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.890 0.940 1.080 1.375 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.430 1.460 1.620 ;
        RECT  1.200 1.430 1.320 1.860 ;
        RECT  0.210 1.740 1.200 1.860 ;
        RECT  0.210 1.005 0.485 1.265 ;
        RECT  0.070 1.005 0.210 1.860 ;
        END
        AntennaGateArea 0.119 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.330 0.570 7.490 2.040 ;
        END
        AntennaDiffArea 0.207 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.090 0.410 7.210 1.935 ;
        RECT  6.745 0.410 7.090 0.530 ;
        RECT  7.055 1.425 7.090 1.935 ;
        RECT  6.760 1.720 7.055 1.840 ;
        RECT  6.500 1.720 6.760 2.100 ;
        RECT  6.575 0.360 6.745 0.530 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.910 1.740 1.170 ;
        END
        AntennaGateArea 0.071 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.225 1.380 3.615 1.620 ;
        RECT  3.105 1.020 3.225 1.620 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.170 -0.210 7.560 0.210 ;
        RECT  6.910 -0.210 7.170 0.290 ;
        RECT  6.050 -0.210 6.910 0.210 ;
        RECT  5.790 -0.210 6.050 0.340 ;
        RECT  4.755 -0.210 5.790 0.210 ;
        RECT  4.495 -0.210 4.755 0.430 ;
        RECT  3.615 -0.210 4.495 0.210 ;
        RECT  3.355 -0.210 3.615 0.420 ;
        RECT  2.950 -0.210 3.355 0.210 ;
        RECT  2.690 -0.210 2.950 0.420 ;
        RECT  1.300 -0.210 2.690 0.210 ;
        RECT  1.040 -0.210 1.300 0.300 ;
        RECT  0.265 -0.210 1.040 0.210 ;
        RECT  0.095 -0.210 0.265 0.495 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.140 2.310 7.560 2.730 ;
        RECT  6.880 2.220 7.140 2.730 ;
        RECT  6.040 2.310 6.880 2.730 ;
        RECT  5.780 1.575 6.040 2.730 ;
        RECT  4.755 2.310 5.780 2.730 ;
        RECT  4.495 2.220 4.755 2.730 ;
        RECT  3.715 2.310 4.495 2.730 ;
        RECT  3.455 2.220 3.715 2.730 ;
        RECT  2.995 2.310 3.455 2.730 ;
        RECT  2.735 2.220 2.995 2.730 ;
        RECT  1.320 2.310 2.735 2.730 ;
        RECT  1.060 2.220 1.320 2.730 ;
        RECT  0.255 2.310 1.060 2.730 ;
        RECT  0.085 1.980 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  6.915 0.650 6.970 1.235 ;
        RECT  6.795 0.650 6.915 1.445 ;
        RECT  6.180 0.650 6.795 0.770 ;
        RECT  6.375 1.325 6.795 1.445 ;
        RECT  6.095 0.975 6.615 1.205 ;
        RECT  6.205 1.325 6.375 1.650 ;
        RECT  5.900 1.325 6.205 1.445 ;
        RECT  5.370 0.975 6.095 1.095 ;
        RECT  5.640 1.215 5.900 1.445 ;
        RECT  5.355 0.370 5.615 0.550 ;
        RECT  5.200 0.705 5.370 1.775 ;
        RECT  5.075 0.430 5.355 0.550 ;
        RECT  5.075 1.980 5.265 2.100 ;
        RECT  4.955 0.430 5.075 2.100 ;
        RECT  4.555 0.620 4.955 0.740 ;
        RECT  2.600 1.980 4.955 2.100 ;
        RECT  4.705 1.000 4.825 1.860 ;
        RECT  3.975 1.740 4.705 1.860 ;
        RECT  4.435 0.620 4.555 1.310 ;
        RECT  4.335 1.050 4.435 1.310 ;
        RECT  4.215 1.495 4.375 1.615 ;
        RECT  4.215 0.330 4.305 0.920 ;
        RECT  4.095 0.330 4.215 1.615 ;
        RECT  3.835 0.330 4.095 0.590 ;
        RECT  3.855 0.755 3.975 1.860 ;
        RECT  3.685 0.755 3.855 0.875 ;
        RECT  2.840 1.740 3.855 1.860 ;
        RECT  3.595 1.000 3.715 1.260 ;
        RECT  3.505 1.000 3.595 1.120 ;
        RECT  3.385 0.540 3.505 1.120 ;
        RECT  2.360 0.540 3.385 0.660 ;
        RECT  2.600 0.780 3.255 0.900 ;
        RECT  2.720 1.260 2.840 1.860 ;
        RECT  2.480 0.780 2.600 2.190 ;
        RECT  2.290 2.020 2.480 2.190 ;
        RECT  2.240 0.540 2.360 1.900 ;
        RECT  2.120 2.020 2.290 2.140 ;
        RECT  2.060 0.540 2.240 0.730 ;
        RECT  2.000 0.920 2.120 2.140 ;
        RECT  1.860 0.920 2.000 1.040 ;
        RECT  1.670 0.380 1.930 0.540 ;
        RECT  1.760 1.660 1.880 2.180 ;
        RECT  0.430 1.980 1.760 2.100 ;
        RECT  0.670 0.420 1.670 0.540 ;
        RECT  0.745 0.660 1.440 0.780 ;
        RECT  0.745 1.500 0.850 1.620 ;
        RECT  0.625 0.660 0.745 1.620 ;
        RECT  0.410 0.380 0.670 0.540 ;
        RECT  0.330 0.660 0.625 0.880 ;
        RECT  0.330 1.455 0.625 1.620 ;
    END
END SDFFX1AD
MACRO SDFFX2AD
    CLASS CORE ;
    FOREIGN SDFFX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.010 1.090 1.375 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.465 1.655 1.610 ;
        RECT  1.440 1.345 1.500 1.610 ;
        RECT  1.240 1.345 1.440 1.800 ;
        RECT  0.210 1.680 1.240 1.800 ;
        RECT  0.210 1.005 0.310 1.265 ;
        RECT  0.090 1.005 0.210 1.800 ;
        END
        AntennaGateArea 0.119 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.330 0.340 7.490 2.020 ;
        END
        AntennaDiffArea 0.373 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.755 1.145 6.930 1.375 ;
        RECT  6.585 0.385 6.755 1.555 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.035 1.890 1.375 ;
        RECT  1.530 1.035 1.750 1.155 ;
        END
        AntennaGateArea 0.071 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.965 1.430 3.430 1.665 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.115 -0.210 7.560 0.210 ;
        RECT  6.945 -0.210 7.115 0.810 ;
        RECT  6.095 -0.210 6.945 0.210 ;
        RECT  5.925 -0.210 6.095 0.440 ;
        RECT  4.750 -0.210 5.925 0.210 ;
        RECT  4.490 -0.210 4.750 0.420 ;
        RECT  3.670 -0.210 4.490 0.210 ;
        RECT  3.475 -0.210 3.670 0.515 ;
        RECT  3.070 -0.210 3.475 0.210 ;
        RECT  2.810 -0.210 3.070 0.540 ;
        RECT  1.280 -0.210 2.810 0.210 ;
        RECT  1.020 -0.210 1.280 0.330 ;
        RECT  0.255 -0.210 1.020 0.210 ;
        RECT  0.085 -0.210 0.255 0.465 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.115 2.310 7.560 2.730 ;
        RECT  6.945 1.995 7.115 2.730 ;
        RECT  6.090 2.310 6.945 2.730 ;
        RECT  5.920 2.005 6.090 2.730 ;
        RECT  4.760 2.310 5.920 2.730 ;
        RECT  4.500 2.255 4.760 2.730 ;
        RECT  3.780 2.310 4.500 2.730 ;
        RECT  3.520 2.220 3.780 2.730 ;
        RECT  3.060 2.310 3.520 2.730 ;
        RECT  2.800 2.220 3.060 2.730 ;
        RECT  1.330 2.310 2.800 2.730 ;
        RECT  1.070 2.220 1.330 2.730 ;
        RECT  0.255 2.310 1.070 2.730 ;
        RECT  0.085 1.940 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  7.090 1.000 7.210 1.840 ;
        RECT  6.415 1.720 7.090 1.840 ;
        RECT  6.295 0.725 6.415 1.840 ;
        RECT  6.245 0.725 6.295 0.895 ;
        RECT  6.245 1.440 6.295 1.840 ;
        RECT  5.800 1.720 6.245 1.840 ;
        RECT  5.725 1.015 6.175 1.275 ;
        RECT  5.680 1.720 5.800 1.980 ;
        RECT  5.340 1.155 5.725 1.275 ;
        RECT  5.100 0.410 5.630 0.530 ;
        RECT  5.460 2.070 5.565 2.190 ;
        RECT  5.305 1.980 5.460 2.190 ;
        RECT  5.220 0.675 5.340 1.650 ;
        RECT  5.100 1.980 5.305 2.100 ;
        RECT  4.980 0.410 5.100 2.100 ;
        RECT  4.620 0.800 4.980 0.920 ;
        RECT  3.375 1.980 4.980 2.100 ;
        RECT  4.740 1.040 4.860 1.860 ;
        RECT  4.020 1.740 4.740 1.860 ;
        RECT  4.500 0.800 4.620 1.255 ;
        RECT  4.380 1.085 4.500 1.255 ;
        RECT  4.260 1.475 4.420 1.595 ;
        RECT  4.300 0.680 4.360 0.940 ;
        RECT  4.260 0.330 4.300 0.940 ;
        RECT  4.140 0.330 4.260 1.595 ;
        RECT  3.950 0.330 4.140 0.450 ;
        RECT  3.900 0.590 4.020 1.860 ;
        RECT  2.640 1.190 3.900 1.310 ;
        RECT  3.790 1.600 3.900 1.860 ;
        RECT  2.370 0.950 3.780 1.070 ;
        RECT  2.610 0.710 3.450 0.830 ;
        RECT  3.175 1.835 3.375 2.100 ;
        RECT  2.560 1.980 3.175 2.100 ;
        RECT  2.490 0.380 2.610 0.830 ;
        RECT  2.300 1.980 2.560 2.135 ;
        RECT  2.130 0.380 2.490 0.500 ;
        RECT  2.250 0.640 2.370 1.845 ;
        RECT  2.130 1.980 2.300 2.100 ;
        RECT  2.010 0.380 2.130 2.100 ;
        RECT  1.770 0.735 2.010 0.855 ;
        RECT  1.755 1.710 1.890 2.085 ;
        RECT  1.695 0.395 1.865 0.615 ;
        RECT  0.440 1.965 1.755 2.085 ;
        RECT  0.605 0.495 1.695 0.615 ;
        RECT  0.560 0.760 1.420 0.880 ;
        RECT  0.560 1.300 0.780 1.560 ;
        RECT  0.435 0.395 0.605 0.615 ;
        RECT  0.440 0.760 0.560 1.560 ;
        RECT  0.330 0.760 0.440 0.880 ;
        RECT  0.330 1.410 0.440 1.560 ;
    END
END SDFFX2AD
MACRO SDFFX4AD
    CLASS CORE ;
    FOREIGN SDFFX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.000 1.080 1.375 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.460 1.470 1.655 1.610 ;
        RECT  1.330 1.430 1.460 1.610 ;
        RECT  1.200 1.430 1.330 1.855 ;
        RECT  0.210 1.735 1.200 1.855 ;
        RECT  0.210 1.005 0.310 1.265 ;
        RECT  0.090 1.005 0.210 1.855 ;
        END
        AntennaGateArea 0.119 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.145 1.005 9.170 1.515 ;
        RECT  9.025 0.400 9.145 2.175 ;
        RECT  8.905 0.400 9.025 0.830 ;
        RECT  8.905 1.485 9.025 2.175 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.185 0.370 8.355 1.545 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.145 1.890 1.375 ;
        RECT  1.570 1.145 1.750 1.350 ;
        END
        AntennaGateArea 0.071 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  2.950 1.430 3.430 1.665 ;
        END
        AntennaGateArea 0.095 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.435 -0.210 9.520 0.210 ;
        RECT  9.265 -0.210 9.435 0.850 ;
        RECT  8.715 -0.210 9.265 0.210 ;
        RECT  8.545 -0.210 8.715 0.820 ;
        RECT  7.995 -0.210 8.545 0.210 ;
        RECT  7.825 -0.210 7.995 0.535 ;
        RECT  7.360 -0.210 7.825 0.210 ;
        RECT  7.100 -0.210 7.360 0.310 ;
        RECT  5.290 -0.210 7.100 0.210 ;
        RECT  5.030 -0.210 5.290 0.670 ;
        RECT  4.180 -0.210 5.030 0.210 ;
        RECT  3.920 -0.210 4.180 0.525 ;
        RECT  3.070 -0.210 3.920 0.210 ;
        RECT  2.810 -0.210 3.070 0.540 ;
        RECT  1.300 -0.210 2.810 0.210 ;
        RECT  1.040 -0.210 1.300 0.375 ;
        RECT  0.265 -0.210 1.040 0.210 ;
        RECT  0.095 -0.210 0.265 0.475 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.435 2.310 9.520 2.730 ;
        RECT  9.265 1.675 9.435 2.730 ;
        RECT  8.715 2.310 9.265 2.730 ;
        RECT  8.545 1.985 8.715 2.730 ;
        RECT  7.995 2.310 8.545 2.730 ;
        RECT  7.825 2.105 7.995 2.730 ;
        RECT  7.490 2.310 7.825 2.730 ;
        RECT  7.230 2.215 7.490 2.730 ;
        RECT  5.490 2.310 7.230 2.730 ;
        RECT  5.230 1.965 5.490 2.730 ;
        RECT  4.790 2.310 5.230 2.730 ;
        RECT  4.530 2.220 4.790 2.730 ;
        RECT  3.780 2.310 4.530 2.730 ;
        RECT  3.520 2.220 3.780 2.730 ;
        RECT  3.060 2.310 3.520 2.730 ;
        RECT  2.800 2.220 3.060 2.730 ;
        RECT  1.320 2.310 2.800 2.730 ;
        RECT  1.060 2.220 1.320 2.730 ;
        RECT  0.255 2.310 1.060 2.730 ;
        RECT  0.085 1.975 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.520 2.520 ;
        LAYER M1 ;
        RECT  8.725 1.015 8.900 1.275 ;
        RECT  8.605 1.015 8.725 1.785 ;
        RECT  8.060 1.665 8.605 1.785 ;
        RECT  7.940 0.685 8.060 1.785 ;
        RECT  7.525 0.685 7.940 0.855 ;
        RECT  7.725 1.665 7.940 1.785 ;
        RECT  7.180 1.030 7.780 1.290 ;
        RECT  7.555 1.410 7.725 2.030 ;
        RECT  6.960 1.910 7.555 2.030 ;
        RECT  7.060 0.620 7.180 1.575 ;
        RECT  6.715 0.620 7.060 0.740 ;
        RECT  6.790 1.405 7.060 1.575 ;
        RECT  6.680 0.900 6.940 1.215 ;
        RECT  6.670 1.405 6.790 2.140 ;
        RECT  6.540 0.380 6.715 0.740 ;
        RECT  6.330 1.095 6.680 1.215 ;
        RECT  6.635 1.405 6.670 1.575 ;
        RECT  6.210 2.020 6.670 2.140 ;
        RECT  6.030 0.380 6.540 0.500 ;
        RECT  6.355 1.695 6.525 1.900 ;
        RECT  5.805 1.695 6.355 1.815 ;
        RECT  6.175 0.670 6.345 0.925 ;
        RECT  6.115 1.095 6.330 1.575 ;
        RECT  5.950 1.965 6.210 2.140 ;
        RECT  5.625 0.805 6.175 0.925 ;
        RECT  5.810 1.375 6.115 1.575 ;
        RECT  5.885 0.380 6.030 0.685 ;
        RECT  5.770 0.565 5.885 0.685 ;
        RECT  4.820 1.455 5.810 1.575 ;
        RECT  5.635 1.695 5.805 2.130 ;
        RECT  5.060 1.695 5.635 1.815 ;
        RECT  5.455 0.670 5.625 0.925 ;
        RECT  4.865 0.805 5.455 0.925 ;
        RECT  4.580 1.210 5.410 1.330 ;
        RECT  4.940 1.695 5.060 2.065 ;
        RECT  4.695 0.675 4.865 0.925 ;
        RECT  4.700 1.455 4.820 2.100 ;
        RECT  4.410 1.980 4.700 2.100 ;
        RECT  4.560 0.355 4.680 0.475 ;
        RECT  4.460 1.210 4.580 1.860 ;
        RECT  4.420 0.355 4.560 0.780 ;
        RECT  4.025 1.740 4.460 1.860 ;
        RECT  4.340 0.660 4.420 0.780 ;
        RECT  4.150 1.980 4.410 2.190 ;
        RECT  4.220 0.660 4.340 1.620 ;
        RECT  3.475 1.980 4.150 2.100 ;
        RECT  3.905 0.675 4.025 1.860 ;
        RECT  3.755 0.675 3.905 0.795 ;
        RECT  3.855 1.190 3.905 1.860 ;
        RECT  2.830 1.190 3.855 1.310 ;
        RECT  2.370 0.950 3.775 1.070 ;
        RECT  3.585 0.625 3.755 0.795 ;
        RECT  3.185 1.885 3.475 2.100 ;
        RECT  2.610 0.710 3.450 0.830 ;
        RECT  2.610 1.980 3.185 2.100 ;
        RECT  2.710 1.190 2.830 1.450 ;
        RECT  2.490 0.385 2.610 0.830 ;
        RECT  2.560 1.980 2.610 2.140 ;
        RECT  2.490 1.980 2.560 2.190 ;
        RECT  2.130 0.385 2.490 0.505 ;
        RECT  2.300 2.020 2.490 2.190 ;
        RECT  2.250 0.640 2.370 1.900 ;
        RECT  2.130 2.020 2.300 2.140 ;
        RECT  2.010 0.385 2.130 2.140 ;
        RECT  1.795 0.890 2.010 1.010 ;
        RECT  1.720 0.495 1.890 0.755 ;
        RECT  1.755 1.780 1.880 2.100 ;
        RECT  0.685 1.980 1.755 2.100 ;
        RECT  0.625 0.495 1.720 0.615 ;
        RECT  1.215 0.760 1.475 1.040 ;
        RECT  0.565 0.760 1.215 0.880 ;
        RECT  0.565 1.480 0.850 1.615 ;
        RECT  0.425 1.980 0.685 2.140 ;
        RECT  0.455 0.395 0.625 0.615 ;
        RECT  0.445 0.760 0.565 1.615 ;
        RECT  0.380 0.760 0.445 0.880 ;
        RECT  0.330 1.480 0.445 1.615 ;
    END
END SDFFX4AD
MACRO SDFFXLAD
    CLASS CORE ;
    FOREIGN SDFFXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.980 1.080 1.240 ;
        RECT  0.910 0.980 1.050 1.435 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.335 1.425 1.460 1.565 ;
        RECT  1.200 1.425 1.335 1.770 ;
        RECT  0.210 1.650 1.200 1.770 ;
        RECT  0.210 1.005 0.485 1.265 ;
        RECT  0.070 1.005 0.210 1.770 ;
        END
        AntennaGateArea 0.119 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.330 0.630 7.490 1.880 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.070 0.470 7.210 1.655 ;
        RECT  6.540 0.470 7.070 0.590 ;
        RECT  6.715 1.535 7.070 1.655 ;
        RECT  6.545 1.535 6.715 1.870 ;
        END
        AntennaDiffArea 0.138 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.420 0.910 1.730 1.180 ;
        END
        AntennaGateArea 0.071 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.225 1.380 3.615 1.620 ;
        RECT  3.105 1.020 3.225 1.620 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.180 -0.210 7.560 0.210 ;
        RECT  6.920 -0.210 7.180 0.330 ;
        RECT  6.015 -0.210 6.920 0.210 ;
        RECT  5.845 -0.210 6.015 0.365 ;
        RECT  4.690 -0.210 5.845 0.210 ;
        RECT  4.690 0.380 4.755 0.500 ;
        RECT  4.570 -0.210 4.690 0.500 ;
        RECT  3.615 -0.210 4.570 0.210 ;
        RECT  4.495 0.380 4.570 0.500 ;
        RECT  3.355 -0.210 3.615 0.420 ;
        RECT  2.950 -0.210 3.355 0.210 ;
        RECT  2.690 -0.210 2.950 0.420 ;
        RECT  1.300 -0.210 2.690 0.210 ;
        RECT  1.040 -0.210 1.300 0.300 ;
        RECT  0.265 -0.210 1.040 0.210 ;
        RECT  0.095 -0.210 0.265 0.495 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.070 2.310 7.560 2.730 ;
        RECT  7.070 1.795 7.140 1.915 ;
        RECT  6.950 1.795 7.070 2.730 ;
        RECT  6.880 1.795 6.950 1.915 ;
        RECT  5.990 2.310 6.950 2.730 ;
        RECT  5.990 1.580 6.060 1.700 ;
        RECT  5.870 1.580 5.990 2.730 ;
        RECT  5.800 1.580 5.870 1.700 ;
        RECT  4.755 2.310 5.870 2.730 ;
        RECT  4.495 2.220 4.755 2.730 ;
        RECT  3.715 2.310 4.495 2.730 ;
        RECT  3.455 2.220 3.715 2.730 ;
        RECT  2.995 2.310 3.455 2.730 ;
        RECT  2.735 2.220 2.995 2.730 ;
        RECT  1.320 2.310 2.735 2.730 ;
        RECT  1.060 2.220 1.320 2.730 ;
        RECT  0.255 2.310 1.060 2.730 ;
        RECT  0.085 1.890 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  6.830 0.710 6.950 1.385 ;
        RECT  6.395 0.710 6.830 0.830 ;
        RECT  6.375 1.265 6.830 1.385 ;
        RECT  6.040 0.950 6.560 1.145 ;
        RECT  6.225 0.625 6.395 0.830 ;
        RECT  6.205 1.265 6.375 1.705 ;
        RECT  5.895 1.265 6.205 1.385 ;
        RECT  5.320 0.950 6.040 1.070 ;
        RECT  5.635 1.190 5.895 1.385 ;
        RECT  5.355 0.370 5.615 0.510 ;
        RECT  5.075 0.390 5.355 0.510 ;
        RECT  5.200 0.650 5.320 1.710 ;
        RECT  5.075 1.905 5.265 2.100 ;
        RECT  4.955 0.390 5.075 2.100 ;
        RECT  4.555 0.620 4.955 0.740 ;
        RECT  2.600 1.980 4.955 2.100 ;
        RECT  4.715 0.980 4.835 1.860 ;
        RECT  3.975 1.740 4.715 1.860 ;
        RECT  4.435 0.620 4.555 1.380 ;
        RECT  4.335 1.120 4.435 1.380 ;
        RECT  4.215 1.500 4.375 1.620 ;
        RECT  4.215 0.460 4.305 0.920 ;
        RECT  4.095 0.330 4.215 1.620 ;
        RECT  3.835 0.330 4.095 0.590 ;
        RECT  3.855 0.755 3.975 1.860 ;
        RECT  3.685 0.755 3.855 0.875 ;
        RECT  2.840 1.740 3.855 1.860 ;
        RECT  3.595 1.000 3.715 1.260 ;
        RECT  3.505 1.000 3.595 1.120 ;
        RECT  3.385 0.540 3.505 1.120 ;
        RECT  2.360 0.540 3.385 0.660 ;
        RECT  2.600 0.780 3.255 0.900 ;
        RECT  2.720 1.260 2.840 1.860 ;
        RECT  2.480 0.780 2.600 2.190 ;
        RECT  2.290 2.020 2.480 2.190 ;
        RECT  2.240 0.540 2.360 1.900 ;
        RECT  2.120 2.020 2.290 2.140 ;
        RECT  2.060 0.540 2.240 0.730 ;
        RECT  2.000 0.850 2.120 2.140 ;
        RECT  1.945 0.850 2.000 1.110 ;
        RECT  1.670 0.380 1.930 0.540 ;
        RECT  1.760 1.710 1.880 2.100 ;
        RECT  0.690 1.980 1.760 2.100 ;
        RECT  0.670 0.420 1.670 0.540 ;
        RECT  0.745 0.660 1.440 0.780 ;
        RECT  0.745 1.270 0.780 1.530 ;
        RECT  0.625 0.660 0.745 1.530 ;
        RECT  0.430 1.890 0.690 2.100 ;
        RECT  0.410 0.380 0.670 0.540 ;
        RECT  0.330 0.660 0.625 0.880 ;
        RECT  0.330 1.410 0.625 1.530 ;
    END
END SDFFXLAD
MACRO SDFFYQX2AD
    CLASS CORE ;
    FOREIGN SDFFYQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.145 1.670 1.335 ;
        RECT  1.200 1.145 1.320 1.405 ;
        RECT  1.145 1.145 1.200 1.335 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 1.470 1.655 1.760 ;
        RECT  0.280 1.640 1.425 1.760 ;
        RECT  0.160 1.015 0.280 1.760 ;
        END
        AntennaGateArea 0.266 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.890 0.410 8.050 2.015 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.945 0.865 2.200 1.260 ;
        END
        AntennaGateArea 0.152 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.670 1.445 4.240 1.610 ;
        END
        AntennaGateArea 0.119 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.585 -0.210 8.120 0.210 ;
        RECT  6.895 -0.210 7.585 0.475 ;
        RECT  5.860 -0.210 6.895 0.210 ;
        RECT  5.600 -0.210 5.860 0.740 ;
        RECT  4.715 -0.210 5.600 0.210 ;
        RECT  4.545 -0.210 4.715 0.750 ;
        RECT  4.020 -0.210 4.545 0.210 ;
        RECT  3.760 -0.210 4.020 0.510 ;
        RECT  1.665 -0.210 3.760 0.210 ;
        RECT  1.405 -0.210 1.665 0.320 ;
        RECT  0.230 -0.210 1.405 0.210 ;
        RECT  0.110 -0.210 0.230 0.860 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.585 2.310 8.120 2.730 ;
        RECT  6.895 2.025 7.585 2.730 ;
        RECT  5.850 2.310 6.895 2.730 ;
        RECT  5.590 2.260 5.850 2.730 ;
        RECT  4.740 2.310 5.590 2.730 ;
        RECT  4.480 2.260 4.740 2.730 ;
        RECT  4.000 2.310 4.480 2.730 ;
        RECT  3.740 2.010 4.000 2.730 ;
        RECT  1.695 2.310 3.740 2.730 ;
        RECT  1.435 2.160 1.695 2.730 ;
        RECT  0.255 2.310 1.435 2.730 ;
        RECT  0.085 1.900 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.120 2.520 ;
        LAYER M1 ;
        RECT  7.650 0.830 7.770 1.695 ;
        RECT  7.360 0.830 7.650 0.950 ;
        RECT  6.870 1.525 7.650 1.695 ;
        RECT  7.110 1.095 7.530 1.215 ;
        RECT  7.240 0.690 7.360 0.950 ;
        RECT  6.990 0.620 7.110 1.215 ;
        RECT  6.410 0.620 6.990 0.740 ;
        RECT  6.750 1.120 6.870 1.695 ;
        RECT  6.410 2.020 6.670 2.190 ;
        RECT  6.340 0.340 6.600 0.500 ;
        RECT  6.290 0.620 6.410 1.730 ;
        RECT  6.145 2.020 6.410 2.140 ;
        RECT  6.100 0.380 6.340 0.500 ;
        RECT  6.220 0.620 6.290 0.740 ;
        RECT  6.100 0.915 6.145 2.140 ;
        RECT  6.025 0.380 6.100 2.140 ;
        RECT  5.980 0.380 6.025 1.035 ;
        RECT  4.315 2.020 6.025 2.140 ;
        RECT  5.665 0.915 5.980 1.035 ;
        RECT  5.785 1.155 5.905 1.900 ;
        RECT  5.065 1.780 5.785 1.900 ;
        RECT  5.545 0.915 5.665 1.390 ;
        RECT  5.430 1.130 5.545 1.390 ;
        RECT  5.290 1.540 5.470 1.660 ;
        RECT  5.350 0.750 5.400 1.010 ;
        RECT  5.290 0.330 5.350 1.010 ;
        RECT  5.170 0.330 5.290 1.660 ;
        RECT  5.090 0.330 5.170 0.450 ;
        RECT  5.050 1.730 5.065 1.900 ;
        RECT  4.930 0.760 5.050 1.900 ;
        RECT  4.860 1.505 4.930 1.900 ;
        RECT  4.480 1.505 4.860 1.625 ;
        RECT  4.600 0.870 4.770 1.355 ;
        RECT  3.250 0.870 4.600 0.990 ;
        RECT  4.360 1.180 4.480 1.625 ;
        RECT  3.480 0.630 4.400 0.750 ;
        RECT  3.590 1.180 4.360 1.300 ;
        RECT  4.195 1.770 4.315 2.140 ;
        RECT  4.145 1.770 4.195 2.090 ;
        RECT  3.200 1.770 4.145 1.890 ;
        RECT  3.360 0.380 3.480 0.750 ;
        RECT  3.250 1.530 3.390 1.650 ;
        RECT  2.625 0.380 3.360 0.500 ;
        RECT  3.200 0.870 3.250 1.650 ;
        RECT  3.080 0.620 3.200 1.650 ;
        RECT  2.940 1.770 3.200 2.190 ;
        RECT  2.745 0.620 3.080 0.740 ;
        RECT  2.885 1.770 2.940 1.890 ;
        RECT  2.765 1.010 2.885 1.890 ;
        RECT  2.625 1.010 2.765 1.130 ;
        RECT  2.505 0.380 2.625 1.130 ;
        RECT  2.345 1.545 2.515 2.000 ;
        RECT  2.340 1.010 2.505 1.130 ;
        RECT  2.240 0.400 2.360 0.660 ;
        RECT  0.885 1.880 2.345 2.000 ;
        RECT  0.930 0.445 2.240 0.565 ;
        RECT  1.440 0.710 1.560 0.970 ;
        RECT  0.660 0.710 1.440 0.830 ;
        RECT  0.660 1.400 0.985 1.520 ;
        RECT  0.715 0.390 0.930 0.565 ;
        RECT  0.715 1.880 0.885 2.155 ;
        RECT  0.670 0.390 0.715 0.510 ;
        RECT  0.540 0.710 0.660 1.520 ;
        RECT  0.400 0.710 0.540 0.880 ;
        RECT  0.400 1.400 0.540 1.520 ;
    END
END SDFFYQX2AD
MACRO SEDFFHQX1AD
    CLASS CORE ;
    FOREIGN SEDFFHQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.100 0.860 1.770 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.390 0.900 3.725 1.020 ;
        RECT  3.270 0.380 3.390 1.020 ;
        RECT  0.820 0.380 3.270 0.500 ;
        RECT  0.700 0.380 0.820 0.560 ;
        RECT  0.505 0.440 0.700 0.560 ;
        RECT  0.350 0.440 0.505 1.480 ;
        RECT  0.330 1.065 0.350 1.480 ;
        END
        AntennaGateArea 0.13 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.520 0.565 11.690 1.945 ;
        END
        AntennaDiffArea 0.21 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.895 1.045 4.015 1.470 ;
        RECT  3.385 1.140 3.895 1.470 ;
        RECT  3.045 1.140 3.385 1.265 ;
        RECT  2.925 1.000 3.045 1.265 ;
        END
        AntennaGateArea 0.1 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.120 2.005 1.455 ;
        END
        AntennaGateArea 0.08 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  5.945 0.920 6.230 1.060 ;
        RECT  5.750 0.920 5.945 1.610 ;
        RECT  5.625 1.190 5.750 1.610 ;
        END
        AntennaGateArea 0.114 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.250 -0.210 11.760 0.210 ;
        RECT  11.130 -0.210 11.250 0.645 ;
        RECT  10.525 -0.210 11.130 0.210 ;
        RECT  10.005 -0.210 10.525 0.260 ;
        RECT  7.610 -0.210 10.005 0.210 ;
        RECT  7.350 -0.210 7.610 0.260 ;
        RECT  6.890 -0.210 7.350 0.210 ;
        RECT  6.630 -0.210 6.890 0.260 ;
        RECT  5.360 -0.210 6.630 0.210 ;
        RECT  5.100 -0.210 5.360 0.260 ;
        RECT  4.275 -0.210 5.100 0.210 ;
        RECT  4.015 -0.210 4.275 0.300 ;
        RECT  3.485 -0.210 4.015 0.210 ;
        RECT  3.225 -0.210 3.485 0.255 ;
        RECT  2.200 -0.210 3.225 0.210 ;
        RECT  1.940 -0.210 2.200 0.260 ;
        RECT  0.580 -0.210 1.940 0.210 ;
        RECT  0.320 -0.210 0.580 0.300 ;
        RECT  0.000 -0.210 0.320 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.350 2.310 11.760 2.730 ;
        RECT  11.090 1.560 11.350 2.730 ;
        RECT  10.430 2.310 11.090 2.730 ;
        RECT  10.260 1.530 10.430 2.730 ;
        RECT  9.055 2.310 10.260 2.730 ;
        RECT  8.795 2.220 9.055 2.730 ;
        RECT  7.495 2.310 8.795 2.730 ;
        RECT  7.235 2.220 7.495 2.730 ;
        RECT  6.885 2.310 7.235 2.730 ;
        RECT  6.625 2.220 6.885 2.730 ;
        RECT  5.790 2.310 6.625 2.730 ;
        RECT  5.530 2.220 5.790 2.730 ;
        RECT  4.375 2.310 5.530 2.730 ;
        RECT  4.115 2.220 4.375 2.730 ;
        RECT  3.695 2.310 4.115 2.730 ;
        RECT  3.435 2.245 3.695 2.730 ;
        RECT  2.915 2.310 3.435 2.730 ;
        RECT  2.655 2.250 2.915 2.730 ;
        RECT  2.490 2.310 2.655 2.730 ;
        RECT  2.230 2.105 2.490 2.730 ;
        RECT  0.580 2.310 2.230 2.730 ;
        RECT  0.320 2.195 0.580 2.730 ;
        RECT  0.000 2.310 0.320 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.760 2.520 ;
        LAYER M1 ;
        RECT  11.185 0.780 11.305 1.410 ;
        RECT  10.890 0.780 11.185 0.900 ;
        RECT  10.860 1.290 11.185 1.410 ;
        RECT  10.625 1.035 11.065 1.155 ;
        RECT  10.770 0.380 10.890 0.900 ;
        RECT  10.690 1.290 10.860 1.785 ;
        RECT  5.265 0.380 10.770 0.500 ;
        RECT  10.385 1.290 10.690 1.410 ;
        RECT  10.505 0.690 10.625 1.155 ;
        RECT  9.835 0.690 10.505 0.810 ;
        RECT  10.265 1.150 10.385 1.410 ;
        RECT  9.955 0.930 10.075 2.190 ;
        RECT  9.735 1.925 9.955 2.190 ;
        RECT  9.715 0.690 9.835 1.740 ;
        RECT  8.525 1.925 9.735 2.045 ;
        RECT  9.615 1.480 9.715 1.740 ;
        RECT  9.475 0.630 9.595 1.260 ;
        RECT  8.095 0.630 9.475 0.750 ;
        RECT  9.355 1.565 9.400 1.780 ;
        RECT  9.230 0.900 9.355 1.780 ;
        RECT  9.095 0.900 9.230 1.020 ;
        RECT  8.845 1.660 9.230 1.780 ;
        RECT  8.990 1.160 9.110 1.420 ;
        RECT  8.385 1.160 8.990 1.280 ;
        RECT  8.585 1.400 8.845 1.780 ;
        RECT  8.440 1.925 8.525 2.190 ;
        RECT  8.265 1.790 8.440 2.190 ;
        RECT  8.310 0.910 8.385 1.280 ;
        RECT  8.310 1.550 8.355 1.670 ;
        RECT  8.170 0.910 8.310 1.670 ;
        RECT  7.975 1.790 8.265 1.910 ;
        RECT  8.125 0.910 8.170 1.030 ;
        RECT  8.095 1.550 8.170 1.670 ;
        RECT  7.755 2.070 8.145 2.190 ;
        RECT  7.970 0.630 8.095 0.780 ;
        RECT  7.855 0.940 7.975 1.910 ;
        RECT  7.320 0.660 7.970 0.780 ;
        RECT  7.515 0.940 7.855 1.060 ;
        RECT  5.505 1.740 7.855 1.860 ;
        RECT  7.635 1.980 7.755 2.190 ;
        RECT  7.450 1.260 7.735 1.430 ;
        RECT  5.150 1.980 7.635 2.100 ;
        RECT  7.320 1.260 7.450 1.620 ;
        RECT  7.200 0.660 7.320 1.620 ;
        RECT  7.070 0.660 7.200 0.780 ;
        RECT  6.240 1.500 7.200 1.620 ;
        RECT  6.670 0.920 7.080 1.180 ;
        RECT  6.530 0.920 6.670 1.380 ;
        RECT  6.410 0.620 6.530 1.380 ;
        RECT  5.905 0.620 6.410 0.740 ;
        RECT  6.120 1.210 6.240 1.620 ;
        RECT  5.505 0.660 5.785 0.780 ;
        RECT  5.385 0.660 5.505 1.860 ;
        RECT  5.145 0.380 5.265 1.550 ;
        RECT  5.025 1.955 5.150 2.100 ;
        RECT  4.905 0.450 5.025 2.100 ;
        RECT  4.625 0.450 4.905 0.575 ;
        RECT  4.890 1.955 4.905 2.100 ;
        RECT  3.850 1.980 4.890 2.100 ;
        RECT  4.665 0.830 4.785 1.860 ;
        RECT  4.595 0.830 4.665 1.000 ;
        RECT  4.610 1.600 4.665 1.860 ;
        RECT  4.505 0.360 4.625 0.620 ;
        RECT  4.475 0.740 4.595 1.000 ;
        RECT  4.330 1.120 4.465 1.715 ;
        RECT  4.210 0.570 4.330 1.715 ;
        RECT  3.615 0.570 4.210 0.740 ;
        RECT  3.975 1.595 4.210 1.715 ;
        RECT  3.730 1.765 3.850 2.100 ;
        RECT  2.970 1.765 3.730 1.885 ;
        RECT  2.730 2.005 3.410 2.125 ;
        RECT  3.115 1.385 3.235 1.645 ;
        RECT  2.790 1.385 3.115 1.505 ;
        RECT  2.850 1.625 2.970 1.885 ;
        RECT  2.790 0.620 2.945 0.740 ;
        RECT  1.870 1.625 2.850 1.745 ;
        RECT  2.670 0.620 2.790 1.505 ;
        RECT  2.610 1.865 2.730 2.125 ;
        RECT  2.365 0.985 2.670 1.245 ;
        RECT  2.110 1.865 2.610 1.985 ;
        RECT  2.245 0.690 2.550 0.810 ;
        RECT  2.245 1.385 2.450 1.505 ;
        RECT  2.125 0.690 2.245 1.505 ;
        RECT  2.030 0.690 2.125 0.810 ;
        RECT  1.990 1.865 2.110 2.140 ;
        RECT  1.910 0.620 2.030 0.810 ;
        RECT  1.100 2.020 1.990 2.140 ;
        RECT  1.390 0.620 1.910 0.740 ;
        RECT  1.750 1.625 1.870 1.900 ;
        RECT  1.630 0.860 1.770 0.980 ;
        RECT  1.150 1.780 1.750 1.900 ;
        RECT  1.510 0.860 1.630 1.630 ;
        RECT  1.350 1.510 1.510 1.630 ;
        RECT  1.270 0.620 1.390 1.210 ;
        RECT  1.030 0.620 1.150 1.900 ;
        RECT  0.840 2.020 1.100 2.180 ;
        RECT  0.720 1.945 0.840 2.180 ;
        RECT  0.230 1.945 0.720 2.065 ;
        RECT  0.210 0.610 0.230 0.870 ;
        RECT  0.210 1.635 0.230 2.065 ;
        RECT  0.090 0.610 0.210 2.065 ;
    END
END SEDFFHQX1AD
MACRO SEDFFHQX2AD
    CLASS CORE ;
    FOREIGN SEDFFHQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.100 0.860 1.770 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.700 0.900 3.895 1.020 ;
        RECT  3.580 0.380 3.700 1.020 ;
        RECT  0.820 0.380 3.580 0.500 ;
        RECT  0.700 0.380 0.820 0.560 ;
        RECT  0.505 0.440 0.700 0.560 ;
        RECT  0.350 0.440 0.505 1.480 ;
        RECT  0.330 1.065 0.350 1.480 ;
        END
        AntennaGateArea 0.128 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.210 0.380 13.370 2.015 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.065 1.005 4.185 1.470 ;
        RECT  3.555 1.140 4.065 1.470 ;
        RECT  3.215 1.140 3.555 1.265 ;
        RECT  3.095 1.000 3.215 1.265 ;
        END
        AntennaGateArea 0.1 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.085 0.860 2.170 1.250 ;
        RECT  1.895 0.860 2.085 1.295 ;
        RECT  1.825 1.175 1.895 1.295 ;
        END
        AntennaGateArea 0.14 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.115 0.920 6.400 1.060 ;
        RECT  5.920 0.920 6.115 1.610 ;
        END
        AntennaGateArea 0.125 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.970 -0.210 13.440 0.210 ;
        RECT  12.850 -0.210 12.970 0.675 ;
        RECT  12.115 -0.210 12.850 0.210 ;
        RECT  11.855 -0.210 12.115 0.260 ;
        RECT  9.855 -0.210 11.855 0.210 ;
        RECT  9.595 -0.210 9.855 0.260 ;
        RECT  9.295 -0.210 9.595 0.210 ;
        RECT  9.035 -0.210 9.295 0.260 ;
        RECT  7.760 -0.210 9.035 0.210 ;
        RECT  7.500 -0.210 7.760 0.260 ;
        RECT  7.030 -0.210 7.500 0.210 ;
        RECT  6.510 -0.210 7.030 0.260 ;
        RECT  5.530 -0.210 6.510 0.210 ;
        RECT  5.270 -0.210 5.530 0.260 ;
        RECT  4.455 -0.210 5.270 0.210 ;
        RECT  4.195 -0.210 4.455 0.330 ;
        RECT  3.655 -0.210 4.195 0.210 ;
        RECT  3.395 -0.210 3.655 0.260 ;
        RECT  2.200 -0.210 3.395 0.210 ;
        RECT  1.940 -0.210 2.200 0.260 ;
        RECT  0.580 -0.210 1.940 0.210 ;
        RECT  0.320 -0.210 0.580 0.300 ;
        RECT  0.000 -0.210 0.320 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.995 2.310 13.440 2.730 ;
        RECT  12.825 1.790 12.995 2.730 ;
        RECT  12.310 2.310 12.825 2.730 ;
        RECT  12.050 1.715 12.310 2.730 ;
        RECT  10.205 2.310 12.050 2.730 ;
        RECT  9.945 2.190 10.205 2.730 ;
        RECT  9.485 2.310 9.945 2.730 ;
        RECT  9.225 2.190 9.485 2.730 ;
        RECT  8.695 2.310 9.225 2.730 ;
        RECT  8.435 2.205 8.695 2.730 ;
        RECT  7.055 2.310 8.435 2.730 ;
        RECT  6.795 2.220 7.055 2.730 ;
        RECT  5.960 2.310 6.795 2.730 ;
        RECT  5.700 2.220 5.960 2.730 ;
        RECT  4.545 2.310 5.700 2.730 ;
        RECT  4.285 2.220 4.545 2.730 ;
        RECT  3.865 2.310 4.285 2.730 ;
        RECT  3.605 2.220 3.865 2.730 ;
        RECT  3.145 2.310 3.605 2.730 ;
        RECT  2.885 2.220 3.145 2.730 ;
        RECT  2.490 2.310 2.885 2.730 ;
        RECT  2.230 2.140 2.490 2.730 ;
        RECT  0.580 2.310 2.230 2.730 ;
        RECT  0.320 2.195 0.580 2.730 ;
        RECT  0.000 2.310 0.320 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 13.440 2.520 ;
        LAYER M1 ;
        RECT  12.920 0.830 13.040 1.595 ;
        RECT  12.570 0.830 12.920 0.950 ;
        RECT  12.090 1.475 12.920 1.595 ;
        RECT  12.330 1.085 12.795 1.255 ;
        RECT  12.450 0.380 12.570 0.950 ;
        RECT  5.435 0.380 12.450 0.500 ;
        RECT  12.210 0.620 12.330 1.255 ;
        RECT  11.205 0.620 12.210 0.740 ;
        RECT  11.970 1.020 12.090 1.595 ;
        RECT  11.730 1.090 11.850 2.140 ;
        RECT  11.585 1.090 11.730 1.210 ;
        RECT  10.445 2.020 11.730 2.140 ;
        RECT  11.490 1.370 11.610 1.660 ;
        RECT  11.465 0.860 11.585 1.210 ;
        RECT  11.205 1.540 11.490 1.660 ;
        RECT  11.325 0.860 11.465 0.980 ;
        RECT  10.685 1.780 11.420 1.900 ;
        RECT  11.085 0.620 11.205 1.660 ;
        RECT  10.750 0.620 11.085 0.740 ;
        RECT  10.805 1.490 11.085 1.660 ;
        RECT  10.620 1.005 10.880 1.265 ;
        RECT  10.565 1.670 10.685 1.900 ;
        RECT  10.500 0.620 10.620 1.265 ;
        RECT  10.335 1.670 10.565 1.790 ;
        RECT  8.045 0.620 10.500 0.740 ;
        RECT  10.325 1.950 10.445 2.140 ;
        RECT  10.335 0.935 10.380 1.055 ;
        RECT  10.215 0.935 10.335 1.790 ;
        RECT  8.275 1.950 10.325 2.070 ;
        RECT  10.120 0.935 10.215 1.055 ;
        RECT  9.335 1.670 10.215 1.790 ;
        RECT  9.845 0.930 9.965 1.550 ;
        RECT  8.795 0.930 9.845 1.050 ;
        RECT  9.215 1.210 9.335 1.790 ;
        RECT  8.795 1.575 8.900 1.745 ;
        RECT  8.675 0.930 8.795 1.745 ;
        RECT  8.365 0.930 8.675 1.050 ;
        RECT  8.020 1.465 8.675 1.585 ;
        RECT  8.045 1.210 8.555 1.330 ;
        RECT  8.195 0.860 8.365 1.050 ;
        RECT  8.155 1.805 8.275 2.070 ;
        RECT  7.730 1.805 8.155 1.925 ;
        RECT  7.925 0.620 8.045 1.330 ;
        RECT  7.850 1.465 8.020 1.685 ;
        RECT  7.490 0.660 7.925 0.780 ;
        RECT  7.470 2.070 7.795 2.190 ;
        RECT  7.730 0.900 7.780 1.160 ;
        RECT  7.610 0.900 7.730 1.925 ;
        RECT  5.675 1.740 7.610 1.860 ;
        RECT  7.370 0.660 7.490 1.620 ;
        RECT  7.350 1.980 7.470 2.190 ;
        RECT  7.240 0.660 7.370 0.780 ;
        RECT  7.350 1.360 7.370 1.620 ;
        RECT  6.410 1.500 7.350 1.620 ;
        RECT  5.195 1.980 7.350 2.100 ;
        RECT  6.840 0.920 7.250 1.180 ;
        RECT  6.700 0.920 6.840 1.380 ;
        RECT  6.580 0.660 6.700 1.380 ;
        RECT  6.335 0.660 6.580 0.780 ;
        RECT  6.290 1.180 6.410 1.620 ;
        RECT  6.075 0.620 6.335 0.780 ;
        RECT  5.675 0.660 5.955 0.780 ;
        RECT  5.555 0.660 5.675 1.860 ;
        RECT  5.315 0.380 5.435 1.550 ;
        RECT  5.075 0.450 5.195 2.100 ;
        RECT  4.820 0.450 5.075 0.575 ;
        RECT  4.020 1.980 5.075 2.100 ;
        RECT  4.835 0.750 4.955 1.860 ;
        RECT  4.620 0.750 4.835 0.920 ;
        RECT  4.755 1.690 4.835 1.860 ;
        RECT  4.650 0.405 4.820 0.575 ;
        RECT  4.500 1.045 4.635 1.715 ;
        RECT  4.380 0.565 4.500 1.715 ;
        RECT  3.860 0.565 4.380 0.735 ;
        RECT  4.145 1.595 4.380 1.715 ;
        RECT  3.900 1.735 4.020 2.100 ;
        RECT  3.140 1.735 3.900 1.855 ;
        RECT  2.860 1.975 3.580 2.095 ;
        RECT  3.260 1.385 3.430 1.590 ;
        RECT  2.960 1.385 3.260 1.505 ;
        RECT  2.980 1.660 3.140 1.855 ;
        RECT  2.960 0.665 3.115 0.785 ;
        RECT  1.870 1.660 2.980 1.780 ;
        RECT  2.840 0.665 2.960 1.505 ;
        RECT  2.740 1.900 2.860 2.095 ;
        RECT  2.755 0.985 2.840 1.245 ;
        RECT  2.110 1.900 2.740 2.020 ;
        RECT  2.635 1.360 2.720 1.530 ;
        RECT  2.515 0.620 2.635 1.530 ;
        RECT  1.390 0.620 2.515 0.740 ;
        RECT  2.210 1.370 2.380 1.540 ;
        RECT  1.630 1.420 2.210 1.540 ;
        RECT  1.990 1.900 2.110 2.140 ;
        RECT  1.100 2.020 1.990 2.140 ;
        RECT  1.750 1.660 1.870 1.900 ;
        RECT  1.630 0.860 1.770 0.980 ;
        RECT  1.150 1.780 1.750 1.900 ;
        RECT  1.510 0.860 1.630 1.660 ;
        RECT  1.340 1.540 1.510 1.660 ;
        RECT  1.270 0.620 1.390 1.210 ;
        RECT  1.030 0.620 1.150 1.900 ;
        RECT  0.840 2.020 1.100 2.190 ;
        RECT  0.720 1.945 0.840 2.190 ;
        RECT  0.230 1.945 0.720 2.065 ;
        RECT  0.210 0.620 0.230 0.880 ;
        RECT  0.210 1.635 0.230 2.065 ;
        RECT  0.090 0.620 0.210 2.065 ;
    END
END SEDFFHQX2AD
MACRO SEDFFHQX4AD
    CLASS CORE ;
    FOREIGN SEDFFHQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.100 0.770 1.655 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.815 0.900 4.185 1.020 ;
        RECT  3.695 0.380 3.815 1.020 ;
        RECT  0.770 0.380 3.695 0.500 ;
        RECT  0.650 0.380 0.770 0.850 ;
        RECT  0.470 0.585 0.650 0.850 ;
        RECT  0.350 0.585 0.470 1.450 ;
        RECT  0.320 1.015 0.350 1.450 ;
        END
        AntennaGateArea 0.128 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.675 1.005 14.790 1.515 ;
        RECT  14.505 0.385 14.675 2.120 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.310 1.000 4.430 1.260 ;
        RECT  3.570 1.140 4.310 1.260 ;
        RECT  3.355 0.865 3.570 1.260 ;
        END
        AntennaGateArea 0.1 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.215 1.120 2.300 1.240 ;
        RECT  1.985 0.910 2.215 1.240 ;
        RECT  1.780 1.120 1.985 1.240 ;
        END
        AntennaGateArea 0.223 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.710 0.910 6.775 1.205 ;
        RECT  6.510 0.765 6.710 1.205 ;
        END
        AntennaGateArea 0.202 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.010 -0.210 15.120 0.210 ;
        RECT  14.890 -0.210 15.010 0.885 ;
        RECT  14.360 -0.210 14.890 0.210 ;
        RECT  14.100 -0.210 14.360 0.500 ;
        RECT  13.385 -0.210 14.100 0.210 ;
        RECT  12.865 -0.210 13.385 0.500 ;
        RECT  10.825 -0.210 12.865 0.210 ;
        RECT  10.565 -0.210 10.825 0.260 ;
        RECT  9.480 -0.210 10.565 0.210 ;
        RECT  8.960 -0.210 9.480 0.260 ;
        RECT  8.130 -0.210 8.960 0.210 ;
        RECT  7.610 -0.210 8.130 0.260 ;
        RECT  6.720 -0.210 7.610 0.210 ;
        RECT  6.460 -0.210 6.720 0.255 ;
        RECT  5.955 -0.210 6.460 0.210 ;
        RECT  5.695 -0.210 5.955 0.260 ;
        RECT  4.670 -0.210 5.695 0.210 ;
        RECT  4.410 -0.210 4.670 0.280 ;
        RECT  3.930 -0.210 4.410 0.210 ;
        RECT  3.670 -0.210 3.930 0.260 ;
        RECT  2.490 -0.210 3.670 0.210 ;
        RECT  1.970 -0.210 2.490 0.260 ;
        RECT  0.530 -0.210 1.970 0.210 ;
        RECT  0.270 -0.210 0.530 0.310 ;
        RECT  0.000 -0.210 0.270 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.010 2.310 15.120 2.730 ;
        RECT  14.890 1.635 15.010 2.730 ;
        RECT  14.315 2.310 14.890 2.730 ;
        RECT  14.145 1.950 14.315 2.730 ;
        RECT  13.790 2.310 14.145 2.730 ;
        RECT  13.620 1.950 13.790 2.730 ;
        RECT  11.200 2.310 13.620 2.730 ;
        RECT  10.940 2.260 11.200 2.730 ;
        RECT  10.420 2.310 10.940 2.730 ;
        RECT  10.160 2.260 10.420 2.730 ;
        RECT  8.115 2.310 10.160 2.730 ;
        RECT  7.595 2.260 8.115 2.730 ;
        RECT  6.100 2.310 7.595 2.730 ;
        RECT  5.840 2.020 6.100 2.730 ;
        RECT  4.900 2.310 5.840 2.730 ;
        RECT  4.640 2.210 4.900 2.730 ;
        RECT  4.120 2.310 4.640 2.730 ;
        RECT  3.860 2.260 4.120 2.730 ;
        RECT  3.340 2.310 3.860 2.730 ;
        RECT  3.080 2.260 3.340 2.730 ;
        RECT  2.760 2.310 3.080 2.730 ;
        RECT  2.240 2.140 2.760 2.730 ;
        RECT  0.590 2.310 2.240 2.730 ;
        RECT  0.330 2.200 0.590 2.730 ;
        RECT  0.000 2.310 0.330 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 15.120 2.520 ;
        LAYER M1 ;
        RECT  14.265 0.620 14.385 1.600 ;
        RECT  13.695 0.620 14.265 0.880 ;
        RECT  13.955 1.430 14.265 1.600 ;
        RECT  13.495 1.050 14.145 1.220 ;
        RECT  13.835 1.430 13.955 1.780 ;
        RECT  13.500 1.660 13.835 1.780 ;
        RECT  12.625 0.620 13.695 0.740 ;
        RECT  13.240 1.660 13.500 2.020 ;
        RECT  13.375 0.860 13.495 1.540 ;
        RECT  12.295 0.860 13.375 0.980 ;
        RECT  12.195 1.420 13.375 1.540 ;
        RECT  11.400 1.140 13.255 1.260 ;
        RECT  9.435 2.020 13.030 2.140 ;
        RECT  11.160 1.745 12.815 1.865 ;
        RECT  12.505 0.380 12.625 0.740 ;
        RECT  5.880 0.380 12.505 0.500 ;
        RECT  12.170 0.620 12.295 0.980 ;
        RECT  11.700 0.620 12.170 0.740 ;
        RECT  11.280 0.660 11.400 1.260 ;
        RECT  7.925 0.660 11.280 0.780 ;
        RECT  10.990 0.955 11.160 1.865 ;
        RECT  10.180 1.745 10.990 1.865 ;
        RECT  10.590 1.000 10.710 1.510 ;
        RECT  9.940 1.000 10.590 1.120 ;
        RECT  10.440 1.390 10.590 1.510 ;
        RECT  10.060 1.305 10.180 1.865 ;
        RECT  9.820 1.000 9.940 1.550 ;
        RECT  9.725 1.430 9.820 1.550 ;
        RECT  9.555 1.430 9.725 1.840 ;
        RECT  8.720 1.430 9.555 1.550 ;
        RECT  9.315 1.685 9.435 2.140 ;
        RECT  8.470 0.965 9.330 1.085 ;
        RECT  8.470 1.685 9.315 1.805 ;
        RECT  9.015 1.930 9.135 2.190 ;
        RECT  6.345 2.020 9.015 2.140 ;
        RECT  8.350 0.965 8.470 1.805 ;
        RECT  7.730 1.685 8.350 1.805 ;
        RECT  7.805 0.660 7.925 1.520 ;
        RECT  7.230 0.660 7.805 0.780 ;
        RECT  7.490 1.400 7.805 1.520 ;
        RECT  7.610 1.685 7.730 1.900 ;
        RECT  7.250 0.965 7.685 1.135 ;
        RECT  6.585 1.780 7.610 1.900 ;
        RECT  7.370 1.400 7.490 1.660 ;
        RECT  6.870 1.540 7.370 1.660 ;
        RECT  7.110 0.965 7.250 1.420 ;
        RECT  6.990 0.640 7.110 1.420 ;
        RECT  6.850 0.640 6.990 0.760 ;
        RECT  6.750 1.400 6.870 1.660 ;
        RECT  6.465 1.495 6.585 1.900 ;
        RECT  6.195 1.495 6.465 1.615 ;
        RECT  6.225 1.735 6.345 2.140 ;
        RECT  6.195 0.640 6.340 0.760 ;
        RECT  5.550 1.735 6.225 1.855 ;
        RECT  6.075 0.640 6.195 1.615 ;
        RECT  5.760 0.380 5.880 1.410 ;
        RECT  5.430 0.570 5.550 2.090 ;
        RECT  5.225 0.570 5.430 0.830 ;
        RECT  4.345 1.970 5.430 2.090 ;
        RECT  5.020 1.140 5.310 1.625 ;
        RECT  4.900 0.520 5.020 1.625 ;
        RECT  4.865 0.520 4.900 0.780 ;
        RECT  4.670 0.920 4.780 1.180 ;
        RECT  4.550 0.590 4.670 1.545 ;
        RECT  4.070 0.590 4.550 0.710 ;
        RECT  4.390 1.425 4.550 1.545 ;
        RECT  4.225 1.780 4.345 2.090 ;
        RECT  3.335 1.780 4.225 1.900 ;
        RECT  3.020 2.020 3.850 2.140 ;
        RECT  3.470 1.385 3.730 1.615 ;
        RECT  3.235 1.385 3.470 1.505 ;
        RECT  3.215 1.660 3.335 1.900 ;
        RECT  3.115 0.620 3.235 1.505 ;
        RECT  1.870 1.660 3.215 1.780 ;
        RECT  3.055 0.620 3.115 1.140 ;
        RECT  3.015 0.880 3.055 1.140 ;
        RECT  2.900 1.900 3.020 2.140 ;
        RECT  2.895 1.280 2.990 1.540 ;
        RECT  2.120 1.900 2.900 2.020 ;
        RECT  2.775 0.620 2.895 1.540 ;
        RECT  1.390 0.620 2.775 0.740 ;
        RECT  1.630 1.420 2.430 1.540 ;
        RECT  2.000 1.900 2.120 2.140 ;
        RECT  1.070 2.020 2.000 2.140 ;
        RECT  1.750 1.660 1.870 1.900 ;
        RECT  1.630 0.860 1.770 0.980 ;
        RECT  1.185 1.780 1.750 1.900 ;
        RECT  1.510 0.860 1.630 1.660 ;
        RECT  1.360 1.510 1.510 1.660 ;
        RECT  1.270 0.620 1.390 1.140 ;
        RECT  1.130 1.020 1.270 1.140 ;
        RECT  1.065 1.600 1.185 1.900 ;
        RECT  1.010 0.620 1.150 0.880 ;
        RECT  0.930 2.020 1.070 2.180 ;
        RECT  1.010 1.600 1.065 1.730 ;
        RECT  0.890 0.620 1.010 1.730 ;
        RECT  0.810 1.900 0.930 2.180 ;
        RECT  0.240 1.900 0.810 2.020 ;
        RECT  0.200 1.610 0.240 2.020 ;
        RECT  0.200 0.600 0.230 0.880 ;
        RECT  0.080 0.600 0.200 2.020 ;
    END
END SEDFFHQX4AD
MACRO SEDFFHQX8AD
    CLASS CORE ;
    FOREIGN SEDFFHQX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.100 0.770 1.655 ;
        END
        AntennaGateArea 0.071 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.780 0.900 6.150 1.020 ;
        RECT  5.660 0.380 5.780 1.020 ;
        RECT  1.370 0.380 5.660 0.500 ;
        RECT  1.110 0.340 1.370 0.500 ;
        RECT  0.770 0.380 1.110 0.500 ;
        RECT  0.650 0.380 0.770 0.850 ;
        RECT  0.470 0.585 0.650 0.850 ;
        RECT  0.350 0.585 0.470 1.450 ;
        RECT  0.320 1.015 0.350 1.450 ;
        END
        AntennaGateArea 0.161 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  18.985 0.370 19.155 2.120 ;
        RECT  18.410 1.005 18.985 1.515 ;
        RECT  18.290 0.340 18.410 2.165 ;
        END
        AntennaDiffArea 0.86 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.275 1.000 6.395 1.260 ;
        RECT  5.535 1.140 6.275 1.260 ;
        RECT  5.320 0.865 5.535 1.260 ;
        END
        AntennaGateArea 0.108 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.825 1.160 3.070 1.330 ;
        RECT  2.550 1.160 2.825 1.280 ;
        END
        AntennaGateArea 0.448 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  8.425 0.910 8.835 1.170 ;
        END
        AntennaGateArea 0.283 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  19.515 -0.210 19.600 0.210 ;
        RECT  19.345 -0.210 19.515 0.800 ;
        RECT  18.795 -0.210 19.345 0.210 ;
        RECT  18.625 -0.210 18.795 0.800 ;
        RECT  18.065 -0.210 18.625 0.210 ;
        RECT  17.895 -0.210 18.065 0.525 ;
        RECT  16.840 -0.210 17.895 0.210 ;
        RECT  16.320 -0.210 16.840 0.255 ;
        RECT  14.125 -0.210 16.320 0.210 ;
        RECT  13.865 -0.210 14.125 0.260 ;
        RECT  13.345 -0.210 13.865 0.210 ;
        RECT  13.085 -0.210 13.345 0.260 ;
        RECT  12.000 -0.210 13.085 0.210 ;
        RECT  11.480 -0.210 12.000 0.260 ;
        RECT  9.935 -0.210 11.480 0.210 ;
        RECT  9.675 -0.210 9.935 0.260 ;
        RECT  8.740 -0.210 9.675 0.210 ;
        RECT  8.480 -0.210 8.740 0.255 ;
        RECT  7.990 -0.210 8.480 0.210 ;
        RECT  7.730 -0.210 7.990 0.260 ;
        RECT  6.635 -0.210 7.730 0.210 ;
        RECT  6.375 -0.210 6.635 0.280 ;
        RECT  5.895 -0.210 6.375 0.210 ;
        RECT  5.635 -0.210 5.895 0.260 ;
        RECT  4.480 -0.210 5.635 0.210 ;
        RECT  3.960 -0.210 4.480 0.230 ;
        RECT  2.950 -0.210 3.960 0.210 ;
        RECT  2.690 -0.210 2.950 0.230 ;
        RECT  0.530 -0.210 2.690 0.210 ;
        RECT  0.270 -0.210 0.530 0.275 ;
        RECT  0.000 -0.210 0.270 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  19.490 2.310 19.600 2.730 ;
        RECT  19.370 1.635 19.490 2.730 ;
        RECT  18.795 2.310 19.370 2.730 ;
        RECT  18.625 1.680 18.795 2.730 ;
        RECT  18.065 2.310 18.625 2.730 ;
        RECT  17.895 1.795 18.065 2.730 ;
        RECT  17.495 2.310 17.895 2.730 ;
        RECT  17.325 1.950 17.495 2.730 ;
        RECT  14.480 2.310 17.325 2.730 ;
        RECT  14.220 2.260 14.480 2.730 ;
        RECT  13.720 2.310 14.220 2.730 ;
        RECT  13.460 2.260 13.720 2.730 ;
        RECT  12.940 2.310 13.460 2.730 ;
        RECT  12.680 2.260 12.940 2.730 ;
        RECT  10.720 2.310 12.680 2.730 ;
        RECT  10.200 2.260 10.720 2.730 ;
        RECT  9.605 2.310 10.200 2.730 ;
        RECT  9.345 2.260 9.605 2.730 ;
        RECT  8.165 2.310 9.345 2.730 ;
        RECT  7.905 2.020 8.165 2.730 ;
        RECT  6.865 2.310 7.905 2.730 ;
        RECT  6.605 2.210 6.865 2.730 ;
        RECT  6.085 2.310 6.605 2.730 ;
        RECT  5.825 2.260 6.085 2.730 ;
        RECT  5.305 2.310 5.825 2.730 ;
        RECT  5.045 2.230 5.305 2.730 ;
        RECT  4.805 2.310 5.045 2.730 ;
        RECT  4.285 2.110 4.805 2.730 ;
        RECT  0.590 2.310 4.285 2.730 ;
        RECT  0.330 2.200 0.590 2.730 ;
        RECT  0.000 2.310 0.330 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 19.600 2.520 ;
        LAYER M1 ;
        RECT  18.045 0.735 18.165 1.600 ;
        RECT  17.570 0.735 18.045 0.880 ;
        RECT  17.635 1.430 18.045 1.600 ;
        RECT  17.040 1.050 17.925 1.220 ;
        RECT  17.515 1.430 17.635 1.780 ;
        RECT  17.405 0.380 17.570 0.880 ;
        RECT  17.110 1.660 17.515 1.780 ;
        RECT  7.945 0.380 17.405 0.500 ;
        RECT  16.990 1.660 17.110 2.090 ;
        RECT  16.920 0.620 17.040 1.540 ;
        RECT  14.605 0.620 16.920 0.740 ;
        RECT  16.615 1.420 16.920 1.540 ;
        RECT  11.955 2.020 16.850 2.140 ;
        RECT  16.655 1.140 16.795 1.260 ;
        RECT  16.535 0.950 16.655 1.260 ;
        RECT  16.610 1.420 16.615 1.850 ;
        RECT  16.440 1.420 16.610 1.900 ;
        RECT  15.515 0.950 16.535 1.070 ;
        RECT  14.960 1.780 16.440 1.900 ;
        RECT  15.250 1.540 16.300 1.660 ;
        RECT  15.130 0.860 15.250 1.660 ;
        RECT  14.435 0.860 15.130 0.980 ;
        RECT  14.815 1.530 15.130 1.660 ;
        RECT  14.195 1.120 14.985 1.240 ;
        RECT  14.645 1.530 14.815 1.800 ;
        RECT  13.955 1.680 14.645 1.800 ;
        RECT  14.315 0.720 14.435 0.980 ;
        RECT  14.075 0.620 14.195 1.240 ;
        RECT  12.875 0.620 14.075 0.740 ;
        RECT  13.835 0.860 13.955 1.800 ;
        RECT  13.465 0.860 13.835 0.980 ;
        RECT  12.700 1.680 13.835 1.800 ;
        RECT  13.210 1.185 13.640 1.355 ;
        RECT  13.090 1.000 13.210 1.355 ;
        RECT  12.460 1.000 13.090 1.120 ;
        RECT  12.615 0.620 12.875 0.780 ;
        RECT  12.580 1.305 12.700 1.800 ;
        RECT  9.990 0.620 12.615 0.740 ;
        RECT  12.340 1.000 12.460 1.550 ;
        RECT  12.245 1.430 12.340 1.550 ;
        RECT  12.075 1.430 12.245 1.840 ;
        RECT  11.455 1.430 12.075 1.550 ;
        RECT  11.835 1.685 11.955 2.140 ;
        RECT  10.990 0.965 11.850 1.085 ;
        RECT  10.990 1.685 11.835 1.805 ;
        RECT  11.535 1.930 11.655 2.190 ;
        RECT  8.410 2.020 11.535 2.140 ;
        RECT  11.285 1.320 11.455 1.550 ;
        RECT  10.870 0.965 10.990 1.805 ;
        RECT  9.995 1.685 10.870 1.805 ;
        RECT  9.875 1.685 9.995 1.900 ;
        RECT  9.870 0.620 9.990 1.520 ;
        RECT  8.650 1.780 9.875 1.900 ;
        RECT  9.290 0.620 9.870 0.780 ;
        RECT  9.555 1.400 9.870 1.520 ;
        RECT  9.315 0.965 9.750 1.135 ;
        RECT  9.435 1.400 9.555 1.660 ;
        RECT  8.935 1.540 9.435 1.660 ;
        RECT  9.170 0.965 9.315 1.420 ;
        RECT  9.055 0.640 9.170 1.420 ;
        RECT  9.005 0.640 9.055 1.135 ;
        RECT  8.910 0.640 9.005 0.760 ;
        RECT  8.815 1.400 8.935 1.660 ;
        RECT  8.530 1.495 8.650 1.900 ;
        RECT  8.260 1.495 8.530 1.615 ;
        RECT  8.260 0.660 8.420 0.780 ;
        RECT  8.290 1.735 8.410 2.140 ;
        RECT  7.615 1.735 8.290 1.855 ;
        RECT  8.140 0.660 8.260 1.615 ;
        RECT  7.825 0.380 7.945 1.410 ;
        RECT  7.525 1.735 7.615 2.090 ;
        RECT  7.395 0.570 7.525 2.090 ;
        RECT  7.170 0.570 7.395 0.830 ;
        RECT  6.310 1.970 7.395 2.090 ;
        RECT  6.985 1.140 7.275 1.625 ;
        RECT  6.865 0.520 6.985 1.625 ;
        RECT  6.830 0.520 6.865 0.780 ;
        RECT  6.635 0.920 6.745 1.180 ;
        RECT  6.515 0.590 6.635 1.545 ;
        RECT  6.035 0.590 6.515 0.710 ;
        RECT  6.355 1.425 6.515 1.545 ;
        RECT  6.190 1.735 6.310 2.090 ;
        RECT  5.300 1.735 6.190 1.855 ;
        RECT  5.785 2.020 5.815 2.140 ;
        RECT  5.555 1.990 5.785 2.140 ;
        RECT  5.435 1.385 5.695 1.615 ;
        RECT  5.045 1.990 5.555 2.110 ;
        RECT  5.200 1.385 5.435 1.505 ;
        RECT  5.180 1.630 5.300 1.855 ;
        RECT  5.080 0.620 5.200 1.505 ;
        RECT  3.705 1.630 5.180 1.750 ;
        RECT  5.020 0.620 5.080 1.120 ;
        RECT  4.925 1.870 5.045 2.110 ;
        RECT  4.980 0.860 5.020 1.120 ;
        RECT  4.860 1.250 4.955 1.510 ;
        RECT  3.950 1.870 4.925 1.990 ;
        RECT  4.860 0.620 4.895 0.740 ;
        RECT  4.740 0.620 4.860 1.510 ;
        RECT  2.160 0.620 4.740 0.740 ;
        RECT  4.450 1.305 4.620 1.510 ;
        RECT  3.455 1.390 4.450 1.510 ;
        RECT  3.830 1.870 3.950 2.140 ;
        RECT  1.120 2.020 3.830 2.140 ;
        RECT  3.585 1.630 3.705 1.900 ;
        RECT  2.030 1.780 3.585 1.900 ;
        RECT  3.335 1.390 3.455 1.630 ;
        RECT  2.400 1.510 3.335 1.630 ;
        RECT  2.400 0.860 3.330 0.980 ;
        RECT  2.280 0.860 2.400 1.630 ;
        RECT  2.130 1.480 2.280 1.630 ;
        RECT  2.040 0.620 2.160 1.110 ;
        RECT  1.540 1.510 2.130 1.630 ;
        RECT  1.810 0.990 2.040 1.110 ;
        RECT  1.770 1.750 2.030 1.900 ;
        RECT  1.750 0.620 1.920 0.790 ;
        RECT  1.200 1.780 1.770 1.900 ;
        RECT  1.010 0.620 1.750 0.740 ;
        RECT  1.540 0.860 1.585 0.980 ;
        RECT  1.410 0.860 1.540 1.630 ;
        RECT  1.325 0.860 1.410 0.980 ;
        RECT  1.080 1.600 1.200 1.900 ;
        RECT  0.860 2.020 1.120 2.180 ;
        RECT  1.010 1.600 1.080 1.730 ;
        RECT  0.890 0.620 1.010 1.730 ;
        RECT  0.840 2.020 0.860 2.140 ;
        RECT  0.720 1.900 0.840 2.140 ;
        RECT  0.240 1.900 0.720 2.020 ;
        RECT  0.200 1.610 0.240 2.020 ;
        RECT  0.200 0.600 0.230 0.880 ;
        RECT  0.080 0.600 0.200 2.020 ;
    END
END SEDFFHQX8AD
MACRO SEDFFTRX1AD
    CLASS CORE ;
    FOREIGN SEDFFTRX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.405 0.865 1.610 1.275 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.040 0.790 1.655 ;
        END
        AntennaGateArea 0.097 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.755 0.235 1.170 ;
        END
        AntennaGateArea 0.057 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.770 1.145 11.970 1.375 ;
        RECT  11.590 0.635 11.770 1.590 ;
        END
        AntennaDiffArea 0.179 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.370 0.645 12.530 1.945 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.145 4.690 1.375 ;
        RECT  4.440 1.145 4.550 1.265 ;
        RECT  4.320 0.945 4.440 1.265 ;
        END
        AntennaGateArea 0.048 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 0.920 3.345 1.180 ;
        RECT  3.150 0.920 3.290 1.375 ;
        END
        AntennaGateArea 0.051 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.230 0.925 6.370 1.380 ;
        RECT  6.150 0.925 6.230 1.185 ;
        END
        AntennaGateArea 0.074 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.155 -0.210 12.600 0.210 ;
        RECT  11.985 -0.210 12.155 0.865 ;
        RECT  11.115 -0.210 11.985 0.210 ;
        RECT  10.855 -0.210 11.115 0.320 ;
        RECT  9.575 -0.210 10.855 0.210 ;
        RECT  9.315 -0.210 9.575 0.415 ;
        RECT  8.425 -0.210 9.315 0.210 ;
        RECT  8.165 -0.210 8.425 0.665 ;
        RECT  7.090 -0.210 8.165 0.210 ;
        RECT  7.065 -0.210 7.090 0.745 ;
        RECT  6.945 -0.210 7.065 0.820 ;
        RECT  6.920 -0.210 6.945 0.745 ;
        RECT  6.500 -0.210 6.920 0.210 ;
        RECT  6.240 -0.210 6.500 0.300 ;
        RECT  4.710 -0.210 6.240 0.210 ;
        RECT  4.450 -0.210 4.710 0.300 ;
        RECT  3.460 -0.210 4.450 0.210 ;
        RECT  3.200 -0.210 3.460 0.300 ;
        RECT  1.440 -0.210 3.200 0.210 ;
        RECT  1.180 -0.210 1.440 0.305 ;
        RECT  0.975 -0.210 1.180 0.210 ;
        RECT  0.805 -0.210 0.975 0.565 ;
        RECT  0.255 -0.210 0.805 0.210 ;
        RECT  0.085 -0.210 0.255 0.555 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.170 2.310 12.600 2.730 ;
        RECT  11.910 1.990 12.170 2.730 ;
        RECT  11.165 2.310 11.910 2.730 ;
        RECT  10.905 2.220 11.165 2.730 ;
        RECT  9.495 2.310 10.905 2.730 ;
        RECT  9.235 2.220 9.495 2.730 ;
        RECT  8.280 2.310 9.235 2.730 ;
        RECT  8.020 2.220 8.280 2.730 ;
        RECT  6.365 2.310 8.020 2.730 ;
        RECT  6.195 2.080 6.365 2.730 ;
        RECT  4.680 2.310 6.195 2.730 ;
        RECT  4.420 2.105 4.680 2.730 ;
        RECT  3.290 2.310 4.420 2.730 ;
        RECT  3.120 1.865 3.290 2.730 ;
        RECT  1.390 2.310 3.120 2.730 ;
        RECT  1.130 2.190 1.390 2.730 ;
        RECT  0.840 2.310 1.130 2.730 ;
        RECT  0.580 2.190 0.840 2.730 ;
        RECT  0.000 2.310 0.580 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 12.600 2.520 ;
        LAYER M1 ;
        RECT  12.130 1.010 12.250 1.870 ;
        RECT  11.470 1.750 12.130 1.870 ;
        RECT  11.350 0.550 11.470 1.870 ;
        RECT  11.280 0.550 11.350 0.720 ;
        RECT  10.815 1.750 11.350 1.870 ;
        RECT  11.030 1.020 11.220 1.280 ;
        RECT  10.910 0.640 11.030 1.280 ;
        RECT  10.230 0.640 10.910 0.760 ;
        RECT  10.695 1.750 10.815 2.140 ;
        RECT  9.695 2.020 10.695 2.140 ;
        RECT  10.425 0.880 10.545 1.900 ;
        RECT  9.925 1.780 10.425 1.900 ;
        RECT  10.060 0.640 10.230 1.635 ;
        RECT  9.830 1.740 9.925 1.900 ;
        RECT  9.795 0.670 9.920 1.620 ;
        RECT  9.360 1.740 9.830 1.860 ;
        RECT  9.750 0.670 9.795 0.840 ;
        RECT  9.635 1.500 9.795 1.620 ;
        RECT  9.600 1.980 9.695 2.140 ;
        RECT  9.610 1.025 9.675 1.285 ;
        RECT  9.490 0.540 9.610 1.285 ;
        RECT  7.855 1.980 9.600 2.100 ;
        RECT  8.715 0.540 9.490 0.660 ;
        RECT  9.240 1.025 9.360 1.860 ;
        RECT  8.955 0.780 9.295 0.900 ;
        RECT  9.210 1.025 9.240 1.285 ;
        RECT  7.615 1.740 9.240 1.860 ;
        RECT  8.955 1.490 9.115 1.610 ;
        RECT  8.835 0.780 8.955 1.610 ;
        RECT  8.620 0.475 8.715 1.300 ;
        RECT  8.595 0.475 8.620 1.575 ;
        RECT  8.450 1.180 8.595 1.575 ;
        RECT  8.150 1.180 8.450 1.300 ;
        RECT  8.325 0.800 8.445 1.060 ;
        RECT  7.740 0.800 8.325 0.920 ;
        RECT  7.890 1.110 8.150 1.300 ;
        RECT  7.735 1.980 7.855 2.140 ;
        RECT  7.620 0.350 7.740 0.920 ;
        RECT  7.060 2.020 7.735 2.140 ;
        RECT  7.570 0.350 7.620 1.620 ;
        RECT  7.300 1.740 7.615 1.900 ;
        RECT  7.500 0.800 7.570 1.620 ;
        RECT  7.420 1.360 7.500 1.620 ;
        RECT  7.300 0.630 7.355 1.155 ;
        RECT  7.235 0.630 7.300 1.900 ;
        RECT  7.180 1.035 7.235 1.900 ;
        RECT  6.660 1.035 7.180 1.155 ;
        RECT  6.940 1.590 7.060 2.140 ;
        RECT  5.770 1.590 6.940 1.710 ;
        RECT  6.700 1.830 6.820 2.135 ;
        RECT  6.015 1.830 6.700 1.950 ;
        RECT  6.540 0.685 6.660 1.155 ;
        RECT  6.090 0.685 6.540 0.805 ;
        RECT  6.010 0.330 6.090 0.805 ;
        RECT  6.010 1.300 6.060 1.470 ;
        RECT  5.895 1.830 6.015 2.140 ;
        RECT  5.890 0.330 6.010 1.470 ;
        RECT  4.960 2.020 5.895 2.140 ;
        RECT  5.830 0.330 5.890 0.450 ;
        RECT  5.650 0.610 5.770 1.900 ;
        RECT  5.460 1.780 5.650 1.900 ;
        RECT  5.380 0.610 5.500 1.660 ;
        RECT  5.290 0.610 5.380 0.870 ;
        RECT  5.315 1.540 5.380 1.660 ;
        RECT  5.185 1.540 5.315 1.875 ;
        RECT  5.170 1.160 5.260 1.420 ;
        RECT  5.145 1.625 5.185 1.875 ;
        RECT  5.070 0.610 5.170 1.420 ;
        RECT  3.915 1.625 5.145 1.745 ;
        RECT  5.050 0.610 5.070 1.495 ;
        RECT  4.950 0.610 5.050 0.780 ;
        RECT  4.810 1.300 5.050 1.495 ;
        RECT  4.840 1.865 4.960 2.140 ;
        RECT  4.830 0.420 4.950 0.780 ;
        RECT  4.810 0.905 4.930 1.180 ;
        RECT  3.540 1.865 4.840 1.985 ;
        RECT  4.160 0.420 4.830 0.540 ;
        RECT  4.680 0.905 4.810 1.025 ;
        RECT  4.560 0.660 4.680 1.025 ;
        RECT  4.155 0.660 4.560 0.780 ;
        RECT  4.155 1.385 4.325 1.505 ;
        RECT  3.990 0.330 4.160 0.540 ;
        RECT  4.035 0.660 4.155 1.505 ;
        RECT  3.990 0.980 4.035 1.240 ;
        RECT  3.870 1.360 3.915 1.745 ;
        RECT  3.750 0.420 3.870 1.745 ;
        RECT  3.080 0.420 3.750 0.540 ;
        RECT  3.505 0.660 3.625 1.505 ;
        RECT  3.420 1.625 3.540 1.985 ;
        RECT  3.320 0.660 3.505 0.780 ;
        RECT  3.410 1.335 3.505 1.505 ;
        RECT  2.785 1.625 3.420 1.745 ;
        RECT  2.985 0.380 3.080 0.540 ;
        RECT  1.970 1.925 3.000 2.045 ;
        RECT  2.480 0.380 2.985 0.500 ;
        RECT  2.865 1.335 2.905 1.505 ;
        RECT  2.695 0.635 2.865 1.505 ;
        RECT  2.665 1.625 2.785 1.805 ;
        RECT  2.450 0.940 2.695 1.060 ;
        RECT  2.230 1.685 2.665 1.805 ;
        RECT  2.375 1.180 2.545 1.565 ;
        RECT  2.330 0.380 2.480 0.710 ;
        RECT  2.330 1.180 2.375 1.300 ;
        RECT  2.325 0.380 2.330 1.300 ;
        RECT  2.210 0.590 2.325 1.300 ;
        RECT  2.110 1.420 2.230 1.805 ;
        RECT  2.090 1.420 2.110 1.540 ;
        RECT  1.970 0.555 2.090 1.540 ;
        RECT  1.850 1.685 1.970 2.045 ;
        RECT  1.730 0.625 1.850 1.565 ;
        RECT  1.120 1.685 1.850 1.805 ;
        RECT  1.530 0.625 1.730 0.745 ;
        RECT  1.645 1.395 1.730 1.565 ;
        RECT  1.550 1.930 1.670 2.190 ;
        RECT  0.485 1.930 1.550 2.050 ;
        RECT  1.000 0.690 1.120 1.805 ;
        RECT  0.870 0.690 1.000 0.950 ;
        RECT  0.485 0.385 0.615 0.840 ;
        RECT  0.445 0.385 0.485 2.050 ;
        RECT  0.365 0.680 0.445 2.050 ;
        RECT  0.085 1.470 0.365 1.640 ;
    END
END SEDFFTRX1AD
MACRO SEDFFTRX2AD
    CLASS CORE ;
    FOREIGN SEDFFTRX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.405 0.865 1.610 1.275 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.040 0.790 1.655 ;
        END
        AntennaGateArea 0.095 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.755 0.235 1.170 ;
        END
        AntennaGateArea 0.055 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.770 1.145 11.970 1.375 ;
        RECT  11.590 0.330 11.770 1.590 ;
        END
        AntennaDiffArea 0.322 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.370 0.330 12.530 2.190 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.145 4.690 1.375 ;
        RECT  4.440 1.145 4.550 1.265 ;
        RECT  4.320 0.945 4.440 1.265 ;
        END
        AntennaGateArea 0.048 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 0.920 3.345 1.180 ;
        RECT  3.150 0.920 3.290 1.375 ;
        END
        AntennaGateArea 0.051 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.230 0.925 6.370 1.380 ;
        RECT  6.150 0.925 6.230 1.185 ;
        END
        AntennaGateArea 0.079 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.155 -0.210 12.600 0.210 ;
        RECT  11.985 -0.210 12.155 0.805 ;
        RECT  11.115 -0.210 11.985 0.210 ;
        RECT  10.855 -0.210 11.115 0.320 ;
        RECT  9.575 -0.210 10.855 0.210 ;
        RECT  9.315 -0.210 9.575 0.415 ;
        RECT  8.425 -0.210 9.315 0.210 ;
        RECT  8.165 -0.210 8.425 0.665 ;
        RECT  7.090 -0.210 8.165 0.210 ;
        RECT  7.065 -0.210 7.090 0.745 ;
        RECT  6.945 -0.210 7.065 0.820 ;
        RECT  6.920 -0.210 6.945 0.745 ;
        RECT  6.500 -0.210 6.920 0.210 ;
        RECT  6.240 -0.210 6.500 0.300 ;
        RECT  4.710 -0.210 6.240 0.210 ;
        RECT  4.450 -0.210 4.710 0.300 ;
        RECT  3.460 -0.210 4.450 0.210 ;
        RECT  3.200 -0.210 3.460 0.300 ;
        RECT  1.440 -0.210 3.200 0.210 ;
        RECT  1.180 -0.210 1.440 0.305 ;
        RECT  0.975 -0.210 1.180 0.210 ;
        RECT  0.805 -0.210 0.975 0.565 ;
        RECT  0.255 -0.210 0.805 0.210 ;
        RECT  0.085 -0.210 0.255 0.565 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.125 2.310 12.600 2.730 ;
        RECT  11.955 1.990 12.125 2.730 ;
        RECT  11.165 2.310 11.955 2.730 ;
        RECT  10.905 2.280 11.165 2.730 ;
        RECT  9.495 2.310 10.905 2.730 ;
        RECT  9.235 2.260 9.495 2.730 ;
        RECT  8.280 2.310 9.235 2.730 ;
        RECT  8.020 2.220 8.280 2.730 ;
        RECT  6.365 2.310 8.020 2.730 ;
        RECT  6.195 2.070 6.365 2.730 ;
        RECT  4.680 2.310 6.195 2.730 ;
        RECT  4.420 2.105 4.680 2.730 ;
        RECT  3.290 2.310 4.420 2.730 ;
        RECT  3.120 1.865 3.290 2.730 ;
        RECT  1.390 2.310 3.120 2.730 ;
        RECT  1.130 2.190 1.390 2.730 ;
        RECT  0.840 2.310 1.130 2.730 ;
        RECT  0.580 2.190 0.840 2.730 ;
        RECT  0.000 2.310 0.580 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 12.600 2.520 ;
        LAYER M1 ;
        RECT  12.130 1.010 12.250 1.870 ;
        RECT  11.470 1.750 12.130 1.870 ;
        RECT  11.350 0.550 11.470 1.870 ;
        RECT  11.280 0.550 11.350 0.720 ;
        RECT  10.815 1.750 11.350 1.870 ;
        RECT  11.030 1.020 11.220 1.280 ;
        RECT  10.910 0.640 11.030 1.280 ;
        RECT  10.280 0.640 10.910 0.760 ;
        RECT  10.695 1.750 10.815 2.140 ;
        RECT  9.180 2.020 10.695 2.140 ;
        RECT  10.425 0.880 10.545 1.900 ;
        RECT  9.420 1.780 10.425 1.900 ;
        RECT  10.110 0.640 10.280 1.635 ;
        RECT  10.065 0.640 10.110 0.760 ;
        RECT  9.795 0.670 9.920 1.660 ;
        RECT  9.750 0.670 9.795 0.840 ;
        RECT  9.635 1.540 9.795 1.660 ;
        RECT  9.610 1.090 9.675 1.350 ;
        RECT  9.490 0.540 9.610 1.350 ;
        RECT  8.715 0.540 9.490 0.660 ;
        RECT  9.360 1.740 9.420 1.900 ;
        RECT  9.300 1.025 9.360 1.900 ;
        RECT  9.240 1.025 9.300 1.860 ;
        RECT  8.955 0.780 9.295 0.900 ;
        RECT  9.210 1.025 9.240 1.285 ;
        RECT  7.615 1.740 9.240 1.860 ;
        RECT  9.090 1.980 9.180 2.140 ;
        RECT  8.955 1.490 9.115 1.610 ;
        RECT  7.855 1.980 9.090 2.100 ;
        RECT  8.835 0.780 8.955 1.610 ;
        RECT  8.620 0.475 8.715 1.300 ;
        RECT  8.595 0.475 8.620 1.575 ;
        RECT  8.450 1.180 8.595 1.575 ;
        RECT  8.150 1.180 8.450 1.300 ;
        RECT  8.325 0.800 8.445 1.060 ;
        RECT  7.740 0.800 8.325 0.920 ;
        RECT  7.890 1.110 8.150 1.300 ;
        RECT  7.735 1.980 7.855 2.140 ;
        RECT  7.620 0.350 7.740 0.920 ;
        RECT  7.060 2.020 7.735 2.140 ;
        RECT  7.570 0.350 7.620 1.620 ;
        RECT  7.300 1.740 7.615 1.900 ;
        RECT  7.500 0.800 7.570 1.620 ;
        RECT  7.420 1.360 7.500 1.620 ;
        RECT  7.300 0.630 7.355 1.155 ;
        RECT  7.235 0.630 7.300 1.900 ;
        RECT  7.180 1.035 7.235 1.900 ;
        RECT  6.660 1.035 7.180 1.155 ;
        RECT  6.940 1.590 7.060 2.140 ;
        RECT  5.770 1.590 6.940 1.710 ;
        RECT  6.700 1.830 6.820 2.135 ;
        RECT  6.015 1.830 6.700 1.950 ;
        RECT  6.540 0.685 6.660 1.155 ;
        RECT  6.090 0.685 6.540 0.805 ;
        RECT  6.010 0.330 6.090 0.805 ;
        RECT  6.010 1.300 6.060 1.470 ;
        RECT  5.895 1.830 6.015 2.140 ;
        RECT  5.890 0.330 6.010 1.470 ;
        RECT  4.960 2.020 5.895 2.140 ;
        RECT  5.830 0.330 5.890 0.450 ;
        RECT  5.650 0.610 5.770 1.900 ;
        RECT  5.460 1.780 5.650 1.900 ;
        RECT  5.380 0.610 5.500 1.660 ;
        RECT  5.290 0.610 5.380 0.870 ;
        RECT  5.315 1.540 5.380 1.660 ;
        RECT  5.185 1.540 5.315 1.875 ;
        RECT  5.170 1.160 5.260 1.420 ;
        RECT  5.145 1.625 5.185 1.875 ;
        RECT  5.070 0.610 5.170 1.420 ;
        RECT  3.915 1.625 5.145 1.745 ;
        RECT  5.050 0.610 5.070 1.495 ;
        RECT  4.950 0.610 5.050 0.780 ;
        RECT  4.810 1.300 5.050 1.495 ;
        RECT  4.840 1.865 4.960 2.140 ;
        RECT  4.830 0.420 4.950 0.780 ;
        RECT  4.810 0.905 4.930 1.180 ;
        RECT  3.540 1.865 4.840 1.985 ;
        RECT  4.160 0.420 4.830 0.540 ;
        RECT  4.680 0.905 4.810 1.025 ;
        RECT  4.560 0.660 4.680 1.025 ;
        RECT  4.155 0.660 4.560 0.780 ;
        RECT  4.155 1.385 4.325 1.505 ;
        RECT  3.990 0.330 4.160 0.540 ;
        RECT  4.035 0.660 4.155 1.505 ;
        RECT  3.990 0.980 4.035 1.240 ;
        RECT  3.870 1.360 3.915 1.745 ;
        RECT  3.750 0.420 3.870 1.745 ;
        RECT  3.080 0.420 3.750 0.540 ;
        RECT  3.505 0.660 3.625 1.505 ;
        RECT  3.420 1.625 3.540 1.985 ;
        RECT  3.320 0.660 3.505 0.780 ;
        RECT  3.410 1.335 3.505 1.505 ;
        RECT  2.785 1.625 3.420 1.745 ;
        RECT  2.985 0.380 3.080 0.540 ;
        RECT  1.970 1.925 3.000 2.045 ;
        RECT  2.480 0.380 2.985 0.500 ;
        RECT  2.865 1.335 2.905 1.505 ;
        RECT  2.695 0.635 2.865 1.505 ;
        RECT  2.665 1.625 2.785 1.805 ;
        RECT  2.450 0.940 2.695 1.060 ;
        RECT  2.230 1.685 2.665 1.805 ;
        RECT  2.375 1.180 2.545 1.565 ;
        RECT  2.330 0.380 2.480 0.710 ;
        RECT  2.330 1.180 2.375 1.300 ;
        RECT  2.325 0.380 2.330 1.300 ;
        RECT  2.210 0.590 2.325 1.300 ;
        RECT  2.110 1.420 2.230 1.805 ;
        RECT  2.090 1.420 2.110 1.540 ;
        RECT  1.970 0.555 2.090 1.540 ;
        RECT  1.850 1.685 1.970 2.045 ;
        RECT  1.730 0.625 1.850 1.565 ;
        RECT  1.120 1.685 1.850 1.805 ;
        RECT  1.530 0.625 1.730 0.745 ;
        RECT  1.645 1.395 1.730 1.565 ;
        RECT  1.550 1.930 1.670 2.190 ;
        RECT  0.485 1.930 1.550 2.050 ;
        RECT  1.000 0.690 1.120 1.805 ;
        RECT  0.870 0.690 1.000 0.950 ;
        RECT  0.485 0.395 0.615 0.840 ;
        RECT  0.445 0.395 0.485 2.050 ;
        RECT  0.365 0.680 0.445 2.050 ;
        RECT  0.085 1.470 0.365 1.640 ;
    END
END SEDFFTRX2AD
MACRO SEDFFTRX4AD
    CLASS CORE ;
    FOREIGN SEDFFTRX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.405 0.865 1.610 1.275 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.055 0.800 1.655 ;
        END
        AntennaGateArea 0.095 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.755 0.235 1.170 ;
        END
        AntennaGateArea 0.055 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.225 0.360 13.395 1.635 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.090 0.360 14.210 1.880 ;
        RECT  14.070 0.360 14.090 2.190 ;
        RECT  13.945 0.360 14.070 0.790 ;
        RECT  13.970 1.410 14.070 2.190 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.145 4.690 1.375 ;
        RECT  4.410 1.145 4.550 1.265 ;
        RECT  4.285 0.995 4.410 1.265 ;
        END
        AntennaGateArea 0.048 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 0.920 3.345 1.180 ;
        RECT  3.150 0.920 3.290 1.375 ;
        END
        AntennaGateArea 0.051 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.230 0.820 6.370 1.380 ;
        RECT  6.120 0.820 6.230 1.080 ;
        END
        AntennaGateArea 0.099 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.475 -0.210 14.560 0.210 ;
        RECT  14.330 -0.210 14.475 0.835 ;
        RECT  13.755 -0.210 14.330 0.210 ;
        RECT  13.585 -0.210 13.755 0.790 ;
        RECT  13.035 -0.210 13.585 0.210 ;
        RECT  12.865 -0.210 13.035 0.500 ;
        RECT  12.320 -0.210 12.865 0.210 ;
        RECT  12.200 -0.210 12.320 0.920 ;
        RECT  10.285 -0.210 12.200 0.210 ;
        RECT  10.025 -0.210 10.285 0.665 ;
        RECT  9.585 -0.210 10.025 0.210 ;
        RECT  9.325 -0.210 9.585 0.415 ;
        RECT  8.420 -0.210 9.325 0.210 ;
        RECT  8.160 -0.210 8.420 0.665 ;
        RECT  7.090 -0.210 8.160 0.210 ;
        RECT  6.920 -0.210 7.090 0.685 ;
        RECT  6.455 -0.210 6.920 0.210 ;
        RECT  6.285 -0.210 6.455 0.255 ;
        RECT  4.705 -0.210 6.285 0.210 ;
        RECT  4.445 -0.210 4.705 0.300 ;
        RECT  3.460 -0.210 4.445 0.210 ;
        RECT  3.200 -0.210 3.460 0.300 ;
        RECT  1.440 -0.210 3.200 0.210 ;
        RECT  1.180 -0.210 1.440 0.305 ;
        RECT  0.975 -0.210 1.180 0.210 ;
        RECT  0.805 -0.210 0.975 0.565 ;
        RECT  0.255 -0.210 0.805 0.210 ;
        RECT  0.085 -0.210 0.255 0.565 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.450 2.310 14.560 2.730 ;
        RECT  14.330 1.410 14.450 2.730 ;
        RECT  13.800 2.310 14.330 2.730 ;
        RECT  13.540 1.995 13.800 2.730 ;
        RECT  13.080 2.310 13.540 2.730 ;
        RECT  12.820 1.995 13.080 2.730 ;
        RECT  12.275 2.310 12.820 2.730 ;
        RECT  12.155 1.660 12.275 2.730 ;
        RECT  10.130 2.310 12.155 2.730 ;
        RECT  9.960 2.265 10.130 2.730 ;
        RECT  9.495 2.310 9.960 2.730 ;
        RECT  9.235 2.220 9.495 2.730 ;
        RECT  8.280 2.310 9.235 2.730 ;
        RECT  8.020 2.220 8.280 2.730 ;
        RECT  6.350 2.310 8.020 2.730 ;
        RECT  6.180 2.115 6.350 2.730 ;
        RECT  4.680 2.310 6.180 2.730 ;
        RECT  4.420 2.105 4.680 2.730 ;
        RECT  3.290 2.310 4.420 2.730 ;
        RECT  3.120 1.885 3.290 2.730 ;
        RECT  1.395 2.310 3.120 2.730 ;
        RECT  1.135 2.190 1.395 2.730 ;
        RECT  0.840 2.310 1.135 2.730 ;
        RECT  0.580 2.190 0.840 2.730 ;
        RECT  0.000 2.310 0.580 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 14.560 2.520 ;
        LAYER M1 ;
        RECT  13.850 1.000 13.940 1.260 ;
        RECT  13.730 1.000 13.850 1.875 ;
        RECT  13.105 1.755 13.730 1.875 ;
        RECT  12.985 0.665 13.105 1.875 ;
        RECT  12.705 0.665 12.985 0.785 ;
        RECT  12.635 1.420 12.985 1.540 ;
        RECT  12.080 1.060 12.865 1.230 ;
        RECT  12.535 0.615 12.705 0.785 ;
        RECT  12.515 1.420 12.635 2.055 ;
        RECT  12.015 1.420 12.515 1.540 ;
        RECT  11.960 0.620 12.080 1.230 ;
        RECT  11.895 1.420 12.015 2.140 ;
        RECT  11.525 0.620 11.960 0.760 ;
        RECT  9.695 2.020 11.895 2.140 ;
        RECT  11.775 0.925 11.830 1.095 ;
        RECT  11.655 0.925 11.775 1.900 ;
        RECT  10.320 1.780 11.655 1.900 ;
        RECT  11.405 0.620 11.525 1.660 ;
        RECT  10.745 0.620 11.405 0.760 ;
        RECT  10.830 1.540 11.405 1.660 ;
        RECT  10.575 0.380 11.365 0.500 ;
        RECT  10.995 1.250 11.255 1.420 ;
        RECT  10.575 1.250 10.995 1.370 ;
        RECT  10.660 1.490 10.830 1.660 ;
        RECT  10.515 0.380 10.575 1.370 ;
        RECT  10.455 0.380 10.515 1.600 ;
        RECT  10.395 0.785 10.455 1.600 ;
        RECT  9.855 0.785 10.395 0.905 ;
        RECT  9.620 1.480 10.395 1.600 ;
        RECT  10.200 1.740 10.320 1.900 ;
        RECT  9.370 1.740 10.200 1.860 ;
        RECT  9.615 1.060 10.120 1.180 ;
        RECT  9.735 0.560 9.855 0.905 ;
        RECT  9.600 1.980 9.695 2.140 ;
        RECT  9.495 0.540 9.615 1.180 ;
        RECT  7.855 1.980 9.600 2.100 ;
        RECT  8.715 0.540 9.495 0.660 ;
        RECT  9.250 1.090 9.370 1.860 ;
        RECT  8.955 0.780 9.285 0.900 ;
        RECT  9.075 1.090 9.250 1.210 ;
        RECT  7.615 1.740 9.250 1.860 ;
        RECT  8.955 1.475 9.115 1.595 ;
        RECT  8.835 0.780 8.955 1.595 ;
        RECT  8.620 0.475 8.715 1.320 ;
        RECT  8.595 0.475 8.620 1.620 ;
        RECT  8.450 1.200 8.595 1.620 ;
        RECT  8.175 1.200 8.450 1.320 ;
        RECT  8.325 0.800 8.445 1.080 ;
        RECT  7.740 0.800 8.325 0.920 ;
        RECT  7.915 1.110 8.175 1.320 ;
        RECT  7.735 1.980 7.855 2.140 ;
        RECT  7.620 0.395 7.740 0.920 ;
        RECT  7.060 2.020 7.735 2.140 ;
        RECT  7.570 0.395 7.620 1.620 ;
        RECT  7.300 1.740 7.615 1.900 ;
        RECT  7.500 0.800 7.570 1.620 ;
        RECT  7.420 1.360 7.500 1.620 ;
        RECT  7.300 0.630 7.355 1.155 ;
        RECT  7.235 0.630 7.300 1.900 ;
        RECT  7.180 1.035 7.235 1.900 ;
        RECT  6.660 1.035 7.180 1.155 ;
        RECT  6.940 1.590 7.060 2.140 ;
        RECT  5.760 1.590 6.940 1.710 ;
        RECT  6.700 1.830 6.820 2.135 ;
        RECT  6.015 1.830 6.700 1.950 ;
        RECT  6.540 0.505 6.660 1.155 ;
        RECT  6.090 0.505 6.540 0.625 ;
        RECT  6.000 0.340 6.090 0.625 ;
        RECT  6.000 1.295 6.060 1.465 ;
        RECT  5.895 1.830 6.015 2.140 ;
        RECT  5.880 0.340 6.000 1.465 ;
        RECT  4.960 2.020 5.895 2.140 ;
        RECT  5.830 0.340 5.880 0.460 ;
        RECT  5.705 0.600 5.760 1.900 ;
        RECT  5.640 0.330 5.705 1.900 ;
        RECT  5.535 0.330 5.640 0.720 ;
        RECT  5.460 1.780 5.640 1.900 ;
        RECT  5.410 0.915 5.500 1.660 ;
        RECT  5.380 0.355 5.410 1.660 ;
        RECT  5.290 0.355 5.380 1.035 ;
        RECT  5.340 1.540 5.380 1.660 ;
        RECT  5.220 1.540 5.340 1.900 ;
        RECT  5.130 0.355 5.290 0.475 ;
        RECT  5.170 1.160 5.260 1.420 ;
        RECT  5.080 1.625 5.220 1.900 ;
        RECT  5.070 0.660 5.170 1.420 ;
        RECT  3.915 1.625 5.080 1.745 ;
        RECT  5.050 0.660 5.070 1.505 ;
        RECT  4.920 0.660 5.050 0.780 ;
        RECT  4.810 1.300 5.050 1.505 ;
        RECT  4.840 1.865 4.960 2.140 ;
        RECT  4.810 0.905 4.930 1.180 ;
        RECT  4.800 0.420 4.920 0.780 ;
        RECT  3.540 1.865 4.840 1.985 ;
        RECT  4.680 0.905 4.810 1.025 ;
        RECT  4.160 0.420 4.800 0.540 ;
        RECT  4.560 0.660 4.680 1.025 ;
        RECT  4.155 0.660 4.560 0.780 ;
        RECT  4.155 1.385 4.330 1.505 ;
        RECT  3.990 0.330 4.160 0.540 ;
        RECT  4.035 0.660 4.155 1.505 ;
        RECT  3.990 0.980 4.035 1.240 ;
        RECT  3.870 1.360 3.915 1.745 ;
        RECT  3.750 0.420 3.870 1.745 ;
        RECT  3.080 0.420 3.750 0.540 ;
        RECT  3.505 0.660 3.625 1.505 ;
        RECT  3.420 1.625 3.540 1.985 ;
        RECT  3.320 0.660 3.505 0.780 ;
        RECT  3.410 1.335 3.505 1.505 ;
        RECT  2.785 1.625 3.420 1.745 ;
        RECT  2.985 0.380 3.080 0.540 ;
        RECT  1.970 1.925 3.000 2.045 ;
        RECT  2.480 0.380 2.985 0.500 ;
        RECT  2.865 1.335 2.905 1.505 ;
        RECT  2.695 0.635 2.865 1.505 ;
        RECT  2.665 1.625 2.785 1.805 ;
        RECT  2.450 0.940 2.695 1.060 ;
        RECT  2.235 1.685 2.665 1.805 ;
        RECT  2.375 1.180 2.545 1.565 ;
        RECT  2.360 0.380 2.480 0.710 ;
        RECT  2.330 1.180 2.375 1.300 ;
        RECT  2.330 0.590 2.360 0.710 ;
        RECT  2.210 0.590 2.330 1.300 ;
        RECT  2.115 1.420 2.235 1.805 ;
        RECT  2.090 1.420 2.115 1.565 ;
        RECT  1.970 0.555 2.090 1.565 ;
        RECT  1.850 1.685 1.970 2.045 ;
        RECT  1.730 0.625 1.850 1.565 ;
        RECT  1.120 1.685 1.850 1.805 ;
        RECT  1.530 0.625 1.730 0.745 ;
        RECT  1.645 1.395 1.730 1.565 ;
        RECT  1.550 1.930 1.670 2.190 ;
        RECT  0.485 1.930 1.550 2.050 ;
        RECT  0.985 0.690 1.120 1.805 ;
        RECT  0.870 0.690 0.985 0.950 ;
        RECT  0.485 0.395 0.615 0.840 ;
        RECT  0.445 0.395 0.485 2.050 ;
        RECT  0.365 0.680 0.445 2.050 ;
        RECT  0.085 1.470 0.365 1.640 ;
    END
END SEDFFTRX4AD
MACRO SEDFFTRXLAD
    CLASS CORE ;
    FOREIGN SEDFFTRXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.405 0.865 1.610 1.275 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.040 0.790 1.655 ;
        END
        AntennaGateArea 0.097 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.755 0.235 1.170 ;
        END
        AntennaGateArea 0.057 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.770 1.145 11.970 1.375 ;
        RECT  11.590 0.645 11.770 1.625 ;
        END
        AntennaDiffArea 0.131 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.370 0.645 12.530 1.685 ;
        END
        AntennaDiffArea 0.143 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.145 4.690 1.375 ;
        RECT  4.440 1.145 4.550 1.265 ;
        RECT  4.320 0.945 4.440 1.265 ;
        END
        AntennaGateArea 0.048 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 0.920 3.345 1.180 ;
        RECT  3.150 0.920 3.290 1.375 ;
        END
        AntennaGateArea 0.051 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.230 0.925 6.370 1.380 ;
        RECT  6.150 0.925 6.230 1.185 ;
        END
        AntennaGateArea 0.074 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.155 -0.210 12.600 0.210 ;
        RECT  11.985 -0.210 12.155 0.860 ;
        RECT  11.115 -0.210 11.985 0.210 ;
        RECT  10.855 -0.210 11.115 0.320 ;
        RECT  9.585 -0.210 10.855 0.210 ;
        RECT  9.325 -0.210 9.585 0.415 ;
        RECT  8.425 -0.210 9.325 0.210 ;
        RECT  8.165 -0.210 8.425 0.665 ;
        RECT  7.090 -0.210 8.165 0.210 ;
        RECT  7.065 -0.210 7.090 0.745 ;
        RECT  6.945 -0.210 7.065 0.820 ;
        RECT  6.920 -0.210 6.945 0.745 ;
        RECT  6.500 -0.210 6.920 0.210 ;
        RECT  6.240 -0.210 6.500 0.300 ;
        RECT  4.710 -0.210 6.240 0.210 ;
        RECT  4.450 -0.210 4.710 0.300 ;
        RECT  3.460 -0.210 4.450 0.210 ;
        RECT  3.200 -0.210 3.460 0.300 ;
        RECT  1.440 -0.210 3.200 0.210 ;
        RECT  1.180 -0.210 1.440 0.305 ;
        RECT  0.975 -0.210 1.180 0.210 ;
        RECT  0.805 -0.210 0.975 0.565 ;
        RECT  0.255 -0.210 0.805 0.210 ;
        RECT  0.085 -0.210 0.255 0.555 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.170 2.310 12.600 2.730 ;
        RECT  11.910 1.990 12.170 2.730 ;
        RECT  11.165 2.310 11.910 2.730 ;
        RECT  10.905 2.220 11.165 2.730 ;
        RECT  9.495 2.310 10.905 2.730 ;
        RECT  9.235 2.220 9.495 2.730 ;
        RECT  8.280 2.310 9.235 2.730 ;
        RECT  8.020 2.220 8.280 2.730 ;
        RECT  6.365 2.310 8.020 2.730 ;
        RECT  6.195 2.080 6.365 2.730 ;
        RECT  4.680 2.310 6.195 2.730 ;
        RECT  4.420 2.105 4.680 2.730 ;
        RECT  3.290 2.310 4.420 2.730 ;
        RECT  3.120 1.865 3.290 2.730 ;
        RECT  1.390 2.310 3.120 2.730 ;
        RECT  1.130 2.190 1.390 2.730 ;
        RECT  0.840 2.310 1.130 2.730 ;
        RECT  0.580 2.190 0.840 2.730 ;
        RECT  0.000 2.310 0.580 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 12.600 2.520 ;
        LAYER M1 ;
        RECT  12.130 1.010 12.250 1.870 ;
        RECT  11.470 1.750 12.130 1.870 ;
        RECT  11.350 0.550 11.470 1.870 ;
        RECT  11.280 0.550 11.350 0.720 ;
        RECT  10.815 1.750 11.350 1.870 ;
        RECT  11.030 1.020 11.220 1.280 ;
        RECT  10.910 0.640 11.030 1.280 ;
        RECT  10.230 0.640 10.910 0.760 ;
        RECT  10.695 1.750 10.815 2.140 ;
        RECT  9.695 2.020 10.695 2.140 ;
        RECT  10.425 0.880 10.545 1.900 ;
        RECT  9.925 1.780 10.425 1.900 ;
        RECT  10.060 0.640 10.230 1.635 ;
        RECT  9.830 1.740 9.925 1.900 ;
        RECT  9.795 0.695 9.920 1.620 ;
        RECT  9.360 1.740 9.830 1.860 ;
        RECT  9.750 0.695 9.795 0.865 ;
        RECT  9.635 1.500 9.795 1.620 ;
        RECT  9.600 1.980 9.695 2.140 ;
        RECT  9.610 1.025 9.675 1.285 ;
        RECT  9.490 0.540 9.610 1.285 ;
        RECT  7.855 1.980 9.600 2.100 ;
        RECT  8.715 0.540 9.490 0.660 ;
        RECT  9.240 1.025 9.360 1.860 ;
        RECT  8.955 0.780 9.295 0.900 ;
        RECT  9.210 1.025 9.240 1.285 ;
        RECT  7.615 1.740 9.240 1.860 ;
        RECT  8.955 1.490 9.115 1.610 ;
        RECT  8.835 0.780 8.955 1.610 ;
        RECT  8.620 0.475 8.715 1.300 ;
        RECT  8.595 0.475 8.620 1.575 ;
        RECT  8.450 1.180 8.595 1.575 ;
        RECT  8.150 1.180 8.450 1.300 ;
        RECT  8.325 0.800 8.445 1.060 ;
        RECT  7.740 0.800 8.325 0.920 ;
        RECT  7.890 1.110 8.150 1.300 ;
        RECT  7.735 1.980 7.855 2.140 ;
        RECT  7.620 0.350 7.740 0.920 ;
        RECT  7.060 2.020 7.735 2.140 ;
        RECT  7.570 0.350 7.620 1.620 ;
        RECT  7.300 1.740 7.615 1.900 ;
        RECT  7.500 0.800 7.570 1.620 ;
        RECT  7.420 1.360 7.500 1.620 ;
        RECT  7.300 0.630 7.355 1.155 ;
        RECT  7.235 0.630 7.300 1.900 ;
        RECT  7.180 1.035 7.235 1.900 ;
        RECT  6.660 1.035 7.180 1.155 ;
        RECT  6.940 1.590 7.060 2.140 ;
        RECT  5.770 1.590 6.940 1.710 ;
        RECT  6.700 1.830 6.820 2.135 ;
        RECT  6.015 1.830 6.700 1.950 ;
        RECT  6.540 0.685 6.660 1.155 ;
        RECT  6.090 0.685 6.540 0.805 ;
        RECT  6.010 0.330 6.090 0.805 ;
        RECT  6.010 1.300 6.060 1.470 ;
        RECT  5.895 1.830 6.015 2.140 ;
        RECT  5.890 0.330 6.010 1.470 ;
        RECT  4.960 2.020 5.895 2.140 ;
        RECT  5.830 0.330 5.890 0.450 ;
        RECT  5.650 0.610 5.770 1.900 ;
        RECT  5.460 1.780 5.650 1.900 ;
        RECT  5.380 0.610 5.500 1.660 ;
        RECT  5.290 0.610 5.380 0.870 ;
        RECT  5.315 1.540 5.380 1.660 ;
        RECT  5.185 1.540 5.315 1.875 ;
        RECT  5.170 1.160 5.260 1.420 ;
        RECT  5.145 1.625 5.185 1.875 ;
        RECT  5.070 0.610 5.170 1.420 ;
        RECT  3.915 1.625 5.145 1.745 ;
        RECT  5.050 0.610 5.070 1.495 ;
        RECT  4.950 0.610 5.050 0.780 ;
        RECT  4.810 1.300 5.050 1.495 ;
        RECT  4.840 1.865 4.960 2.140 ;
        RECT  4.830 0.420 4.950 0.780 ;
        RECT  4.810 0.905 4.930 1.180 ;
        RECT  3.540 1.865 4.840 1.985 ;
        RECT  4.160 0.420 4.830 0.540 ;
        RECT  4.680 0.905 4.810 1.025 ;
        RECT  4.560 0.660 4.680 1.025 ;
        RECT  4.155 0.660 4.560 0.780 ;
        RECT  4.155 1.385 4.325 1.505 ;
        RECT  3.990 0.330 4.160 0.540 ;
        RECT  4.035 0.660 4.155 1.505 ;
        RECT  3.990 0.980 4.035 1.240 ;
        RECT  3.870 1.360 3.915 1.745 ;
        RECT  3.750 0.420 3.870 1.745 ;
        RECT  3.080 0.420 3.750 0.540 ;
        RECT  3.505 0.660 3.625 1.505 ;
        RECT  3.420 1.625 3.540 1.985 ;
        RECT  3.320 0.660 3.505 0.780 ;
        RECT  3.410 1.335 3.505 1.505 ;
        RECT  2.785 1.625 3.420 1.745 ;
        RECT  2.985 0.380 3.080 0.540 ;
        RECT  1.970 1.925 3.000 2.045 ;
        RECT  2.480 0.380 2.985 0.500 ;
        RECT  2.865 1.335 2.905 1.505 ;
        RECT  2.695 0.635 2.865 1.505 ;
        RECT  2.665 1.625 2.785 1.805 ;
        RECT  2.450 0.940 2.695 1.060 ;
        RECT  2.230 1.685 2.665 1.805 ;
        RECT  2.375 1.180 2.545 1.565 ;
        RECT  2.330 0.380 2.480 0.710 ;
        RECT  2.330 1.180 2.375 1.300 ;
        RECT  2.325 0.380 2.330 1.300 ;
        RECT  2.210 0.590 2.325 1.300 ;
        RECT  2.110 1.420 2.230 1.805 ;
        RECT  2.090 1.420 2.110 1.540 ;
        RECT  1.970 0.555 2.090 1.540 ;
        RECT  1.850 1.685 1.970 2.045 ;
        RECT  1.730 0.625 1.850 1.565 ;
        RECT  1.120 1.685 1.850 1.805 ;
        RECT  1.530 0.625 1.730 0.745 ;
        RECT  1.645 1.395 1.730 1.565 ;
        RECT  1.550 1.930 1.670 2.190 ;
        RECT  0.485 1.930 1.550 2.050 ;
        RECT  1.000 0.690 1.120 1.805 ;
        RECT  0.870 0.690 1.000 0.950 ;
        RECT  0.485 0.385 0.615 0.840 ;
        RECT  0.445 0.385 0.485 2.050 ;
        RECT  0.365 0.680 0.445 2.050 ;
        RECT  0.085 1.470 0.365 1.640 ;
    END
END SEDFFTRXLAD
MACRO SEDFFX1AD
    CLASS CORE ;
    FOREIGN SEDFFX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.580 0.910 1.935 1.090 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.915 1.120 1.095 ;
        RECT  0.600 0.865 1.050 1.095 ;
        END
        AntennaGateArea 0.088 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.850 1.425 8.890 1.920 ;
        RECT  8.730 0.625 8.850 1.920 ;
        END
        AntennaDiffArea 0.207 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.250 0.865 8.370 1.860 ;
        RECT  8.130 0.865 8.250 1.095 ;
        RECT  7.660 1.740 8.250 1.860 ;
        RECT  8.010 0.605 8.130 1.095 ;
        END
        AntennaDiffArea 0.183 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.750 0.535 1.890 ;
        RECT  0.110 1.750 0.370 2.140 ;
        END
        AntennaGateArea 0.088 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 0.910 2.495 1.290 ;
        END
        AntennaGateArea 0.04 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.500 1.130 4.855 1.355 ;
        END
        AntennaGateArea 0.077 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.560 -0.210 8.960 0.210 ;
        RECT  8.300 -0.210 8.560 0.745 ;
        RECT  7.540 -0.210 8.300 0.210 ;
        RECT  7.280 -0.210 7.540 0.445 ;
        RECT  6.085 -0.210 7.280 0.210 ;
        RECT  5.825 -0.210 6.085 0.415 ;
        RECT  4.870 -0.210 5.825 0.210 ;
        RECT  4.610 -0.210 4.870 0.415 ;
        RECT  1.730 -0.210 4.610 0.210 ;
        RECT  1.470 -0.210 1.730 0.505 ;
        RECT  0.590 -0.210 1.470 0.210 ;
        RECT  0.330 -0.210 0.590 0.300 ;
        RECT  0.000 -0.210 0.330 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.540 2.310 8.960 2.730 ;
        RECT  8.280 2.220 8.540 2.730 ;
        RECT  7.540 2.310 8.280 2.730 ;
        RECT  7.280 2.220 7.540 2.730 ;
        RECT  6.290 2.310 7.280 2.730 ;
        RECT  6.030 2.220 6.290 2.730 ;
        RECT  5.180 2.310 6.030 2.730 ;
        RECT  4.920 2.220 5.180 2.730 ;
        RECT  4.460 2.310 4.920 2.730 ;
        RECT  4.200 2.220 4.460 2.730 ;
        RECT  1.400 2.310 4.200 2.730 ;
        RECT  1.140 2.060 1.400 2.730 ;
        RECT  0.610 2.310 1.140 2.730 ;
        RECT  0.490 2.010 0.610 2.730 ;
        RECT  0.000 2.310 0.490 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.960 2.520 ;
        LAYER M1 ;
        RECT  8.490 1.005 8.610 2.100 ;
        RECT  7.300 1.980 8.490 2.100 ;
        RECT  8.010 1.330 8.130 1.590 ;
        RECT  7.890 1.330 8.010 1.450 ;
        RECT  7.770 0.755 7.890 1.450 ;
        RECT  7.570 0.755 7.770 0.875 ;
        RECT  7.300 1.330 7.770 1.450 ;
        RECT  7.480 1.000 7.650 1.210 ;
        RECT  7.040 1.000 7.480 1.120 ;
        RECT  7.180 1.300 7.300 2.100 ;
        RECT  3.975 1.980 7.180 2.100 ;
        RECT  6.920 0.755 7.040 1.800 ;
        RECT  6.760 0.375 7.020 0.570 ;
        RECT  6.690 0.755 6.920 1.015 ;
        RECT  6.660 1.680 6.920 1.800 ;
        RECT  6.570 1.385 6.800 1.520 ;
        RECT  6.570 0.450 6.760 0.570 ;
        RECT  6.450 0.450 6.570 1.520 ;
        RECT  6.150 1.085 6.450 1.205 ;
        RECT  6.205 0.375 6.325 0.655 ;
        RECT  5.420 0.535 6.205 0.655 ;
        RECT  6.030 1.085 6.150 1.860 ;
        RECT  5.910 1.085 6.030 1.345 ;
        RECT  4.000 1.740 6.030 1.860 ;
        RECT  5.780 1.500 5.910 1.620 ;
        RECT  5.650 0.810 5.780 1.620 ;
        RECT  5.610 0.810 5.650 1.320 ;
        RECT  5.540 1.060 5.610 1.320 ;
        RECT  5.420 1.500 5.530 1.620 ;
        RECT  5.300 0.535 5.420 1.620 ;
        RECT  5.215 0.535 5.300 0.995 ;
        RECT  4.380 1.500 5.300 1.620 ;
        RECT  5.095 1.120 5.180 1.380 ;
        RECT  5.060 0.620 5.095 1.380 ;
        RECT  4.975 0.620 5.060 1.340 ;
        RECT  3.980 0.620 4.975 0.740 ;
        RECT  4.430 0.860 4.690 1.005 ;
        RECT  4.000 0.860 4.430 0.980 ;
        RECT  4.260 1.360 4.380 1.620 ;
        RECT  3.880 0.860 4.000 1.860 ;
        RECT  3.860 0.475 3.980 0.740 ;
        RECT  3.855 1.980 3.975 2.140 ;
        RECT  3.670 0.860 3.880 0.980 ;
        RECT  3.405 0.620 3.860 0.740 ;
        RECT  3.300 2.020 3.855 2.140 ;
        RECT  3.640 1.120 3.760 1.900 ;
        RECT  2.140 0.380 3.670 0.500 ;
        RECT  3.405 1.120 3.640 1.240 ;
        RECT  1.850 1.750 3.450 1.870 ;
        RECT  3.285 0.620 3.405 1.240 ;
        RECT  3.040 2.020 3.300 2.180 ;
        RECT  2.810 0.930 3.160 1.050 ;
        RECT  1.295 0.625 3.040 0.745 ;
        RECT  1.640 2.020 2.820 2.140 ;
        RECT  2.690 0.930 2.810 1.630 ;
        RECT  2.420 1.470 2.690 1.630 ;
        RECT  0.230 1.510 2.420 1.630 ;
        RECT  1.420 1.270 2.070 1.390 ;
        RECT  1.520 1.820 1.640 2.140 ;
        RECT  0.760 1.820 1.520 1.940 ;
        RECT  1.300 0.875 1.420 1.390 ;
        RECT  0.480 1.270 1.300 1.390 ;
        RECT  1.125 0.540 1.295 0.745 ;
        RECT  0.480 0.620 0.980 0.740 ;
        RECT  0.360 0.620 0.480 1.390 ;
        RECT  0.110 0.550 0.230 1.630 ;
    END
END SEDFFX1AD
MACRO SEDFFX2AD
    CLASS CORE ;
    FOREIGN SEDFFX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.865 2.135 1.095 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.600 0.865 1.150 1.095 ;
        END
        AntennaGateArea 0.129 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.130 1.425 9.170 2.190 ;
        RECT  9.010 0.330 9.130 2.190 ;
        END
        AntennaDiffArea 0.373 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.530 0.865 8.650 1.860 ;
        RECT  8.410 0.865 8.530 1.095 ;
        RECT  7.940 1.740 8.530 1.860 ;
        RECT  8.290 0.330 8.410 1.095 ;
        END
        AntennaDiffArea 0.349 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.750 0.535 1.890 ;
        RECT  0.110 1.750 0.370 2.140 ;
        END
        AntennaGateArea 0.122 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 0.860 2.555 1.135 ;
        END
        AntennaGateArea 0.075 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.780 1.130 5.135 1.355 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.840 -0.210 9.240 0.210 ;
        RECT  8.580 -0.210 8.840 0.745 ;
        RECT  7.775 -0.210 8.580 0.210 ;
        RECT  7.605 -0.210 7.775 0.400 ;
        RECT  6.270 -0.210 7.605 0.210 ;
        RECT  6.010 -0.210 6.270 0.415 ;
        RECT  5.150 -0.210 6.010 0.210 ;
        RECT  4.890 -0.210 5.150 0.415 ;
        RECT  1.940 -0.210 4.890 0.210 ;
        RECT  1.680 -0.210 1.940 0.450 ;
        RECT  0.630 -0.210 1.680 0.210 ;
        RECT  0.370 -0.210 0.630 0.300 ;
        RECT  0.000 -0.210 0.370 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.770 2.310 9.240 2.730 ;
        RECT  8.510 2.220 8.770 2.730 ;
        RECT  7.770 2.310 8.510 2.730 ;
        RECT  7.510 2.220 7.770 2.730 ;
        RECT  6.570 2.310 7.510 2.730 ;
        RECT  6.310 2.220 6.570 2.730 ;
        RECT  5.460 2.310 6.310 2.730 ;
        RECT  5.200 2.220 5.460 2.730 ;
        RECT  4.830 2.310 5.200 2.730 ;
        RECT  4.570 2.265 4.830 2.730 ;
        RECT  1.680 2.310 4.570 2.730 ;
        RECT  1.420 2.065 1.680 2.730 ;
        RECT  0.610 2.310 1.420 2.730 ;
        RECT  0.490 2.010 0.610 2.730 ;
        RECT  0.000 2.310 0.490 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.240 2.520 ;
        LAYER M1 ;
        RECT  8.770 1.005 8.890 2.100 ;
        RECT  7.580 1.980 8.770 2.100 ;
        RECT  8.290 1.330 8.410 1.590 ;
        RECT  8.170 1.330 8.290 1.450 ;
        RECT  8.050 0.755 8.170 1.450 ;
        RECT  7.850 0.755 8.050 0.875 ;
        RECT  7.580 1.330 8.050 1.450 ;
        RECT  7.760 1.000 7.930 1.210 ;
        RECT  7.320 1.000 7.760 1.120 ;
        RECT  7.460 1.300 7.580 2.100 ;
        RECT  4.305 1.980 7.460 2.100 ;
        RECT  7.190 0.350 7.330 0.470 ;
        RECT  7.200 0.825 7.320 1.800 ;
        RECT  6.945 0.825 7.200 0.995 ;
        RECT  6.940 1.680 7.200 1.800 ;
        RECT  7.070 0.350 7.190 0.705 ;
        RECT  6.825 1.400 7.080 1.520 ;
        RECT  6.825 0.585 7.070 0.705 ;
        RECT  6.705 0.585 6.825 1.520 ;
        RECT  6.430 1.085 6.705 1.205 ;
        RECT  6.515 0.330 6.655 0.450 ;
        RECT  6.395 0.330 6.515 0.655 ;
        RECT  6.310 1.085 6.430 1.860 ;
        RECT  5.700 0.535 6.395 0.655 ;
        RECT  6.190 1.085 6.310 1.345 ;
        RECT  4.290 1.740 6.310 1.860 ;
        RECT  6.060 1.500 6.190 1.620 ;
        RECT  5.930 0.810 6.060 1.620 ;
        RECT  5.890 0.810 5.930 1.320 ;
        RECT  5.820 1.060 5.890 1.320 ;
        RECT  5.700 1.500 5.810 1.620 ;
        RECT  5.580 0.535 5.700 1.620 ;
        RECT  5.495 0.535 5.580 0.995 ;
        RECT  4.660 1.500 5.580 1.620 ;
        RECT  5.375 1.120 5.460 1.380 ;
        RECT  5.255 0.620 5.375 1.380 ;
        RECT  4.260 0.620 5.255 0.740 ;
        RECT  4.710 0.860 4.970 1.005 ;
        RECT  4.290 0.860 4.710 0.980 ;
        RECT  4.540 1.360 4.660 1.620 ;
        RECT  4.185 1.980 4.305 2.140 ;
        RECT  4.170 0.860 4.290 1.860 ;
        RECT  4.140 0.475 4.260 0.740 ;
        RECT  3.570 2.020 4.185 2.140 ;
        RECT  3.950 0.860 4.170 0.980 ;
        RECT  3.685 0.620 4.140 0.740 ;
        RECT  3.930 1.120 4.050 1.900 ;
        RECT  2.420 0.380 3.950 0.500 ;
        RECT  3.685 1.120 3.930 1.240 ;
        RECT  2.130 1.750 3.730 1.870 ;
        RECT  3.565 0.620 3.685 1.240 ;
        RECT  3.310 2.020 3.570 2.190 ;
        RECT  2.800 0.900 3.440 1.020 ;
        RECT  1.970 0.620 3.320 0.740 ;
        RECT  1.920 2.020 3.100 2.140 ;
        RECT  2.680 0.900 2.800 1.630 ;
        RECT  0.230 1.510 2.680 1.630 ;
        RECT  1.550 1.270 2.200 1.390 ;
        RECT  1.850 0.570 1.970 0.740 ;
        RECT  1.800 1.820 1.920 2.140 ;
        RECT  1.490 0.570 1.850 0.690 ;
        RECT  1.040 1.820 1.800 1.940 ;
        RECT  1.430 0.810 1.550 1.390 ;
        RECT  1.320 0.505 1.490 0.690 ;
        RECT  0.480 1.270 1.430 1.390 ;
        RECT  0.480 0.620 1.010 0.740 ;
        RECT  0.360 0.620 0.480 1.390 ;
        RECT  0.110 0.550 0.230 1.630 ;
    END
END SEDFFX2AD
MACRO SEDFFX4AD
    CLASS CORE ;
    FOREIGN SEDFFX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.575 0.865 1.975 1.085 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 0.865 1.075 1.095 ;
        END
        AntennaGateArea 0.129 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.035 0.355 11.130 1.920 ;
        RECT  10.990 0.355 11.035 2.180 ;
        RECT  10.865 0.355 10.990 0.785 ;
        RECT  10.865 1.490 10.990 2.180 ;
        END
        AntennaDiffArea 0.422 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.145 0.355 10.315 1.635 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.750 0.535 1.910 ;
        END
        AntennaGateArea 0.126 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.205 0.910 2.555 1.140 ;
        END
        AntennaGateArea 0.078 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.785 1.130 5.135 1.355 ;
        END
        AntennaGateArea 0.09 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.395 -0.210 11.480 0.210 ;
        RECT  11.250 -0.210 11.395 0.830 ;
        RECT  10.675 -0.210 11.250 0.210 ;
        RECT  10.505 -0.210 10.675 0.785 ;
        RECT  9.955 -0.210 10.505 0.210 ;
        RECT  9.785 -0.210 9.955 0.575 ;
        RECT  9.175 -0.210 9.785 0.210 ;
        RECT  8.915 -0.210 9.175 0.310 ;
        RECT  7.855 -0.210 8.915 0.210 ;
        RECT  7.595 -0.210 7.855 0.310 ;
        RECT  6.555 -0.210 7.595 0.210 ;
        RECT  6.295 -0.210 6.555 0.500 ;
        RECT  5.270 -0.210 6.295 0.210 ;
        RECT  4.750 -0.210 5.270 0.415 ;
        RECT  1.760 -0.210 4.750 0.210 ;
        RECT  1.500 -0.210 1.760 0.500 ;
        RECT  0.600 -0.210 1.500 0.210 ;
        RECT  0.340 -0.210 0.600 0.300 ;
        RECT  0.000 -0.210 0.340 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.390 2.310 11.480 2.730 ;
        RECT  11.250 1.445 11.390 2.730 ;
        RECT  10.675 2.310 11.250 2.730 ;
        RECT  10.505 1.995 10.675 2.730 ;
        RECT  10.000 2.310 10.505 2.730 ;
        RECT  9.740 1.995 10.000 2.730 ;
        RECT  9.350 2.310 9.740 2.730 ;
        RECT  9.090 2.220 9.350 2.730 ;
        RECT  7.960 2.310 9.090 2.730 ;
        RECT  7.700 2.220 7.960 2.730 ;
        RECT  6.700 2.310 7.700 2.730 ;
        RECT  6.440 2.220 6.700 2.730 ;
        RECT  5.460 2.310 6.440 2.730 ;
        RECT  5.200 2.220 5.460 2.730 ;
        RECT  4.670 2.310 5.200 2.730 ;
        RECT  4.410 2.220 4.670 2.730 ;
        RECT  1.650 2.310 4.410 2.730 ;
        RECT  1.390 1.990 1.650 2.730 ;
        RECT  0.555 2.310 1.390 2.730 ;
        RECT  0.385 2.035 0.555 2.730 ;
        RECT  0.000 2.310 0.385 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.480 2.520 ;
        LAYER M1 ;
        RECT  10.660 1.020 10.860 1.280 ;
        RECT  10.540 1.020 10.660 1.875 ;
        RECT  10.025 1.755 10.540 1.875 ;
        RECT  9.905 0.695 10.025 1.875 ;
        RECT  9.525 0.695 9.905 0.815 ;
        RECT  9.530 1.400 9.905 1.520 ;
        RECT  9.050 1.080 9.785 1.210 ;
        RECT  9.410 1.400 9.530 2.100 ;
        RECT  9.355 0.525 9.525 0.815 ;
        RECT  4.300 1.980 9.410 2.100 ;
        RECT  8.930 0.430 9.050 1.850 ;
        RECT  7.205 0.430 8.930 0.550 ;
        RECT  7.070 1.730 8.930 1.850 ;
        RECT  8.690 0.670 8.810 1.610 ;
        RECT  8.265 0.670 8.690 0.790 ;
        RECT  8.450 0.910 8.570 1.560 ;
        RECT  7.345 1.440 8.450 1.560 ;
        RECT  8.145 0.670 8.265 1.315 ;
        RECT  7.605 1.195 8.145 1.315 ;
        RECT  7.845 0.950 7.985 1.070 ;
        RECT  7.725 0.670 7.845 1.070 ;
        RECT  6.725 0.670 7.725 0.790 ;
        RECT  7.485 0.910 7.605 1.315 ;
        RECT  6.965 0.910 7.485 1.030 ;
        RECT  7.215 1.200 7.345 1.610 ;
        RECT  6.695 1.490 7.215 1.610 ;
        RECT  6.945 0.380 7.205 0.550 ;
        RECT  6.845 0.910 6.965 1.370 ;
        RECT  6.290 1.250 6.845 1.370 ;
        RECT  6.465 0.620 6.725 1.105 ;
        RECT  6.575 1.490 6.695 1.860 ;
        RECT  4.370 1.740 6.575 1.860 ;
        RECT  5.705 0.620 6.465 0.740 ;
        RECT  6.030 1.250 6.290 1.620 ;
        RECT  5.945 0.860 6.175 0.980 ;
        RECT  5.945 1.250 6.030 1.370 ;
        RECT  5.825 0.860 5.945 1.370 ;
        RECT  5.705 1.500 5.770 1.620 ;
        RECT  5.585 0.620 5.705 1.620 ;
        RECT  5.495 0.620 5.585 0.995 ;
        RECT  4.620 1.500 5.585 1.620 ;
        RECT  5.375 1.120 5.465 1.380 ;
        RECT  5.255 0.545 5.375 1.380 ;
        RECT  4.260 0.545 5.255 0.665 ;
        RECT  4.370 0.860 4.960 1.005 ;
        RECT  4.500 1.360 4.620 1.620 ;
        RECT  4.250 0.860 4.370 1.860 ;
        RECT  4.180 1.980 4.300 2.140 ;
        RECT  4.140 0.460 4.260 0.740 ;
        RECT  3.950 0.860 4.250 1.005 ;
        RECT  4.090 1.360 4.250 1.620 ;
        RECT  3.580 2.020 4.180 2.140 ;
        RECT  3.825 0.620 4.140 0.740 ;
        RECT  3.915 1.750 4.130 1.870 ;
        RECT  2.200 0.380 3.950 0.500 ;
        RECT  3.825 1.160 3.915 1.870 ;
        RECT  3.795 0.620 3.825 1.870 ;
        RECT  3.705 0.620 3.795 1.280 ;
        RECT  3.555 1.610 3.675 1.870 ;
        RECT  3.320 2.020 3.580 2.190 ;
        RECT  2.115 1.750 3.555 1.870 ;
        RECT  3.280 0.760 3.400 1.125 ;
        RECT  2.930 1.005 3.280 1.125 ;
        RECT  1.335 0.620 3.160 0.740 ;
        RECT  1.920 1.990 3.100 2.110 ;
        RECT  2.810 1.005 2.930 1.630 ;
        RECT  2.670 1.175 2.810 1.630 ;
        RECT  0.230 1.510 2.670 1.630 ;
        RECT  1.455 1.270 2.210 1.390 ;
        RECT  1.800 1.750 1.920 2.110 ;
        RECT  1.010 1.750 1.800 1.870 ;
        RECT  1.285 0.885 1.455 1.390 ;
        RECT  1.165 0.540 1.335 0.740 ;
        RECT  0.470 1.270 1.285 1.390 ;
        RECT  0.470 0.620 0.980 0.740 ;
        RECT  0.350 0.620 0.470 1.390 ;
        RECT  0.110 0.550 0.230 1.630 ;
    END
END SEDFFX4AD
MACRO SEDFFXLAD
    CLASS CORE ;
    FOREIGN SEDFFXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.580 0.910 1.935 1.090 ;
        END
        AntennaGateArea 0.04 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.915 1.120 1.095 ;
        RECT  0.600 0.865 1.050 1.095 ;
        END
        AntennaGateArea 0.088 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.450 0.680 8.610 1.690 ;
        END
        AntennaDiffArea 0.143 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.910 0.760 8.050 1.645 ;
        RECT  7.600 0.760 7.910 0.880 ;
        RECT  7.735 1.475 7.910 1.645 ;
        END
        AntennaDiffArea 0.143 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.750 0.535 1.890 ;
        RECT  0.110 1.750 0.370 2.140 ;
        END
        AntennaGateArea 0.088 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 0.910 2.495 1.290 ;
        END
        AntennaGateArea 0.04 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.500 1.130 4.855 1.355 ;
        END
        AntennaGateArea 0.076 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.250 -0.210 8.680 0.210 ;
        RECT  7.990 -0.210 8.250 0.400 ;
        RECT  7.405 -0.210 7.990 0.210 ;
        RECT  7.235 -0.210 7.405 0.365 ;
        RECT  6.085 -0.210 7.235 0.210 ;
        RECT  5.825 -0.210 6.085 0.415 ;
        RECT  4.870 -0.210 5.825 0.210 ;
        RECT  4.610 -0.210 4.870 0.415 ;
        RECT  1.730 -0.210 4.610 0.210 ;
        RECT  1.470 -0.210 1.730 0.505 ;
        RECT  0.590 -0.210 1.470 0.210 ;
        RECT  0.330 -0.210 0.590 0.300 ;
        RECT  0.000 -0.210 0.330 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.285 2.310 8.680 2.730 ;
        RECT  8.115 2.005 8.285 2.730 ;
        RECT  7.520 2.310 8.115 2.730 ;
        RECT  7.260 2.220 7.520 2.730 ;
        RECT  6.290 2.310 7.260 2.730 ;
        RECT  6.030 2.220 6.290 2.730 ;
        RECT  5.180 2.310 6.030 2.730 ;
        RECT  4.920 2.220 5.180 2.730 ;
        RECT  4.460 2.310 4.920 2.730 ;
        RECT  4.200 2.220 4.460 2.730 ;
        RECT  1.400 2.310 4.200 2.730 ;
        RECT  1.140 2.060 1.400 2.730 ;
        RECT  0.610 2.310 1.140 2.730 ;
        RECT  0.490 2.010 0.610 2.730 ;
        RECT  0.000 2.310 0.490 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.680 2.520 ;
        LAYER M1 ;
        RECT  8.210 0.520 8.330 1.885 ;
        RECT  7.830 0.520 8.210 0.640 ;
        RECT  7.980 1.765 8.210 1.885 ;
        RECT  7.860 1.765 7.980 2.100 ;
        RECT  7.300 1.980 7.860 2.100 ;
        RECT  7.570 0.400 7.830 0.640 ;
        RECT  7.490 1.000 7.610 1.535 ;
        RECT  7.040 1.000 7.490 1.120 ;
        RECT  7.180 1.300 7.300 2.100 ;
        RECT  3.975 1.980 7.180 2.100 ;
        RECT  6.920 0.755 7.040 1.800 ;
        RECT  6.760 0.375 7.020 0.570 ;
        RECT  6.690 0.755 6.920 1.015 ;
        RECT  6.660 1.680 6.920 1.800 ;
        RECT  6.570 1.385 6.800 1.520 ;
        RECT  6.570 0.450 6.760 0.570 ;
        RECT  6.450 0.450 6.570 1.520 ;
        RECT  6.150 1.085 6.450 1.205 ;
        RECT  6.205 0.430 6.325 0.690 ;
        RECT  5.420 0.570 6.205 0.690 ;
        RECT  6.030 1.085 6.150 1.860 ;
        RECT  5.910 1.085 6.030 1.345 ;
        RECT  4.000 1.740 6.030 1.860 ;
        RECT  5.780 1.500 5.910 1.620 ;
        RECT  5.650 0.810 5.780 1.620 ;
        RECT  5.610 0.810 5.650 1.320 ;
        RECT  5.540 1.060 5.610 1.320 ;
        RECT  5.420 1.500 5.530 1.620 ;
        RECT  5.300 0.570 5.420 1.620 ;
        RECT  5.215 0.570 5.300 0.995 ;
        RECT  4.380 1.500 5.300 1.620 ;
        RECT  5.095 1.120 5.180 1.380 ;
        RECT  5.060 0.620 5.095 1.380 ;
        RECT  4.975 0.620 5.060 1.340 ;
        RECT  3.980 0.620 4.975 0.740 ;
        RECT  4.430 0.860 4.690 1.005 ;
        RECT  4.000 0.860 4.430 0.980 ;
        RECT  4.260 1.360 4.380 1.620 ;
        RECT  3.880 0.860 4.000 1.860 ;
        RECT  3.860 0.475 3.980 0.740 ;
        RECT  3.855 1.980 3.975 2.140 ;
        RECT  3.670 0.860 3.880 0.980 ;
        RECT  3.405 0.620 3.860 0.740 ;
        RECT  3.300 2.020 3.855 2.140 ;
        RECT  3.640 1.120 3.760 1.900 ;
        RECT  2.140 0.380 3.670 0.500 ;
        RECT  3.405 1.120 3.640 1.240 ;
        RECT  1.850 1.750 3.450 1.870 ;
        RECT  3.285 0.620 3.405 1.240 ;
        RECT  3.040 2.020 3.300 2.180 ;
        RECT  2.810 0.930 3.160 1.050 ;
        RECT  1.295 0.625 3.040 0.745 ;
        RECT  1.640 2.020 2.820 2.140 ;
        RECT  2.690 0.930 2.810 1.630 ;
        RECT  2.420 1.470 2.690 1.630 ;
        RECT  0.230 1.510 2.420 1.630 ;
        RECT  1.420 1.270 2.070 1.390 ;
        RECT  1.520 1.820 1.640 2.140 ;
        RECT  0.760 1.820 1.520 1.940 ;
        RECT  1.300 0.875 1.420 1.390 ;
        RECT  0.480 1.270 1.300 1.390 ;
        RECT  1.125 0.540 1.295 0.745 ;
        RECT  0.480 0.620 0.980 0.740 ;
        RECT  0.360 0.620 0.480 1.390 ;
        RECT  0.110 0.550 0.230 1.630 ;
    END
END SEDFFXLAD
MACRO SMDFFHQX1AD
    CLASS CORE ;
    FOREIGN SMDFFHQX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.335 0.780 1.655 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.490 0.910 3.820 1.030 ;
        RECT  3.370 0.680 3.490 1.030 ;
        RECT  3.260 0.680 3.370 0.800 ;
        RECT  3.140 0.380 3.260 0.800 ;
        RECT  0.770 0.380 3.140 0.500 ;
        RECT  0.650 0.380 0.770 1.200 ;
        RECT  0.340 0.865 0.650 1.200 ;
        END
        AntennaGateArea 0.128 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.970 1.020 4.175 1.330 ;
        RECT  3.645 1.160 3.970 1.330 ;
        RECT  3.100 1.160 3.645 1.280 ;
        RECT  2.980 1.020 3.100 1.280 ;
        END
        AntennaGateArea 0.1 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.960 0.635 11.130 1.915 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.980 0.910 2.215 1.375 ;
        RECT  1.760 1.115 1.980 1.375 ;
        END
        AntennaGateArea 0.05 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 0.865 5.530 1.375 ;
        END
        AntennaGateArea 0.05 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  5.905 0.840 6.425 1.050 ;
        END
        AntennaGateArea 0.114 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.735 -0.210 11.200 0.210 ;
        RECT  10.565 -0.210 10.735 0.300 ;
        RECT  10.265 -0.210 10.565 0.210 ;
        RECT  10.095 -0.210 10.265 0.300 ;
        RECT  8.665 -0.210 10.095 0.210 ;
        RECT  8.495 -0.210 8.665 0.255 ;
        RECT  7.410 -0.210 8.495 0.210 ;
        RECT  7.240 -0.210 7.410 0.255 ;
        RECT  6.330 -0.210 7.240 0.210 ;
        RECT  6.160 -0.210 6.330 0.255 ;
        RECT  5.780 -0.210 6.160 0.210 ;
        RECT  5.610 -0.210 5.780 0.365 ;
        RECT  4.290 -0.210 5.610 0.210 ;
        RECT  4.120 -0.210 4.290 0.415 ;
        RECT  3.595 -0.210 4.120 0.210 ;
        RECT  3.425 -0.210 3.595 0.305 ;
        RECT  2.165 -0.210 3.425 0.210 ;
        RECT  1.995 -0.210 2.165 0.255 ;
        RECT  0.530 -0.210 1.995 0.210 ;
        RECT  0.360 -0.210 0.530 0.340 ;
        RECT  0.000 -0.210 0.360 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.755 2.310 11.200 2.730 ;
        RECT  10.585 1.455 10.755 2.730 ;
        RECT  10.075 2.310 10.585 2.730 ;
        RECT  9.905 1.715 10.075 2.730 ;
        RECT  8.795 2.310 9.905 2.730 ;
        RECT  8.625 2.245 8.795 2.730 ;
        RECT  7.135 2.310 8.625 2.730 ;
        RECT  6.965 2.240 7.135 2.730 ;
        RECT  5.725 2.310 6.965 2.730 ;
        RECT  5.555 2.240 5.725 2.730 ;
        RECT  4.265 2.310 5.555 2.730 ;
        RECT  4.095 2.240 4.265 2.730 ;
        RECT  3.665 2.310 4.095 2.730 ;
        RECT  3.495 2.240 3.665 2.730 ;
        RECT  3.025 2.310 3.495 2.730 ;
        RECT  2.855 2.235 3.025 2.730 ;
        RECT  1.565 2.310 2.855 2.730 ;
        RECT  1.395 2.235 1.565 2.730 ;
        RECT  0.540 2.310 1.395 2.730 ;
        RECT  0.370 2.195 0.540 2.730 ;
        RECT  0.000 2.310 0.370 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.200 2.520 ;
        LAYER M1 ;
        RECT  10.580 1.020 10.840 1.280 ;
        RECT  10.460 0.420 10.580 1.280 ;
        RECT  9.520 0.420 10.460 0.540 ;
        RECT  10.325 1.375 10.375 1.545 ;
        RECT  10.155 0.735 10.325 1.545 ;
        RECT  9.890 1.020 10.155 1.280 ;
        RECT  9.640 0.660 9.760 2.125 ;
        RECT  9.630 2.005 9.640 2.125 ;
        RECT  9.110 2.005 9.630 2.170 ;
        RECT  9.420 0.420 9.520 0.860 ;
        RECT  9.400 0.420 9.420 1.590 ;
        RECT  9.260 0.660 9.400 1.590 ;
        RECT  9.020 0.330 9.280 0.500 ;
        RECT  8.200 2.005 9.110 2.125 ;
        RECT  8.980 0.700 9.100 1.880 ;
        RECT  8.295 0.380 9.020 0.500 ;
        RECT  8.840 0.700 8.980 0.820 ;
        RECT  8.915 1.410 8.980 1.880 ;
        RECT  8.320 1.760 8.915 1.880 ;
        RECT  8.605 0.980 8.860 1.240 ;
        RECT  8.415 0.730 8.605 1.580 ;
        RECT  8.085 0.730 8.415 0.850 ;
        RECT  7.570 1.460 8.415 1.580 ;
        RECT  8.015 0.340 8.295 0.500 ;
        RECT  7.595 1.095 8.210 1.265 ;
        RECT  8.080 1.740 8.200 2.125 ;
        RECT  7.825 0.640 8.085 0.850 ;
        RECT  7.450 1.740 8.080 1.860 ;
        RECT  7.210 0.380 8.015 0.500 ;
        RECT  5.015 2.000 7.950 2.120 ;
        RECT  7.450 0.840 7.595 1.265 ;
        RECT  7.330 0.840 7.450 1.860 ;
        RECT  5.770 1.740 7.330 1.860 ;
        RECT  7.090 0.380 7.210 1.580 ;
        RECT  6.900 0.380 7.090 0.755 ;
        RECT  6.800 1.410 7.090 1.580 ;
        RECT  6.760 0.910 6.870 1.290 ;
        RECT  6.540 1.410 6.800 1.620 ;
        RECT  6.565 0.510 6.760 1.290 ;
        RECT  6.150 1.170 6.565 1.290 ;
        RECT  6.270 1.410 6.540 1.580 ;
        RECT  5.890 1.170 6.150 1.440 ;
        RECT  5.770 0.540 6.085 0.700 ;
        RECT  5.650 0.540 5.770 1.860 ;
        RECT  5.270 1.495 5.415 1.705 ;
        RECT  5.270 0.555 5.400 0.725 ;
        RECT  5.140 0.555 5.270 1.705 ;
        RECT  4.895 0.510 5.015 2.120 ;
        RECT  4.840 1.400 4.895 2.120 ;
        RECT  3.750 2.000 4.840 2.120 ;
        RECT  4.720 1.020 4.775 1.280 ;
        RECT  4.600 0.540 4.720 1.855 ;
        RECT  4.535 0.540 4.600 0.800 ;
        RECT  4.455 1.735 4.600 1.855 ;
        RECT  4.415 1.020 4.475 1.280 ;
        RECT  4.295 0.560 4.415 1.605 ;
        RECT  3.680 0.560 4.295 0.730 ;
        RECT  4.050 1.485 4.295 1.605 ;
        RECT  3.630 1.640 3.750 2.120 ;
        RECT  2.880 1.640 3.630 1.760 ;
        RECT  3.240 1.880 3.500 2.100 ;
        RECT  2.800 1.400 3.380 1.520 ;
        RECT  1.150 1.980 3.240 2.100 ;
        RECT  2.800 0.660 2.990 0.780 ;
        RECT  2.695 1.640 2.880 1.860 ;
        RECT  2.680 0.660 2.800 1.520 ;
        RECT  1.225 1.740 2.695 1.860 ;
        RECT  2.390 0.620 2.560 1.545 ;
        RECT  2.300 0.620 2.390 0.780 ;
        RECT  1.400 0.620 2.300 0.740 ;
        RECT  1.640 1.500 2.020 1.620 ;
        RECT  1.640 0.860 1.780 0.980 ;
        RECT  1.520 0.860 1.640 1.620 ;
        RECT  1.280 0.620 1.400 1.520 ;
        RECT  1.160 1.690 1.225 1.860 ;
        RECT  1.040 0.680 1.160 1.860 ;
        RECT  0.780 1.980 1.150 2.165 ;
        RECT  0.660 1.790 0.780 2.165 ;
        RECT  0.255 1.790 0.660 1.910 ;
        RECT  0.205 0.595 0.255 0.770 ;
        RECT  0.205 1.730 0.255 1.910 ;
        RECT  0.085 0.595 0.205 1.910 ;
    END
END SMDFFHQX1AD
MACRO SMDFFHQX2AD
    CLASS CORE ;
    FOREIGN SMDFFHQX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.260 0.880 1.610 ;
        RECT  0.585 1.470 0.630 1.610 ;
        END
        AntennaGateArea 0.048 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.500 0.925 3.935 1.045 ;
        RECT  3.380 0.590 3.500 1.045 ;
        RECT  3.310 0.590 3.380 0.710 ;
        RECT  3.190 0.380 3.310 0.710 ;
        RECT  0.910 0.380 3.190 0.500 ;
        RECT  0.790 0.380 0.910 1.140 ;
        RECT  0.490 1.020 0.790 1.140 ;
        RECT  0.430 1.020 0.490 1.375 ;
        RECT  0.310 1.020 0.430 1.540 ;
        END
        AntennaGateArea 0.128 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.075 1.010 4.195 1.330 ;
        RECT  3.945 1.165 4.075 1.330 ;
        RECT  3.205 1.165 3.945 1.285 ;
        RECT  3.085 0.940 3.205 1.285 ;
        END
        AntennaGateArea 0.1 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.810 0.350 11.970 2.170 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 1.070 2.175 1.375 ;
        END
        AntennaGateArea 0.077 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.635 0.820 5.810 1.375 ;
        RECT  5.535 0.820 5.635 1.080 ;
        END
        AntennaGateArea 0.077 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.185 0.830 6.505 1.050 ;
        END
        AntennaGateArea 0.117 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.525 -0.210 12.040 0.210 ;
        RECT  11.355 -0.210 11.525 0.305 ;
        RECT  10.790 -0.210 11.355 0.210 ;
        RECT  10.620 -0.210 10.790 0.305 ;
        RECT  8.985 -0.210 10.620 0.210 ;
        RECT  8.725 -0.210 8.985 0.280 ;
        RECT  7.470 -0.210 8.725 0.210 ;
        RECT  7.300 -0.210 7.470 0.415 ;
        RECT  6.370 -0.210 7.300 0.210 ;
        RECT  5.650 -0.210 6.370 0.290 ;
        RECT  4.310 -0.210 5.650 0.210 ;
        RECT  3.530 -0.210 4.310 0.335 ;
        RECT  2.165 -0.210 3.530 0.210 ;
        RECT  1.995 -0.210 2.165 0.255 ;
        RECT  0.575 -0.210 1.995 0.210 ;
        RECT  0.405 -0.210 0.575 0.475 ;
        RECT  0.000 -0.210 0.405 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.595 2.310 12.040 2.730 ;
        RECT  11.425 1.400 11.595 2.730 ;
        RECT  11.160 2.310 11.425 2.730 ;
        RECT  10.990 1.900 11.160 2.730 ;
        RECT  9.450 2.310 10.990 2.730 ;
        RECT  9.280 2.260 9.450 2.730 ;
        RECT  8.870 2.310 9.280 2.730 ;
        RECT  8.700 2.260 8.870 2.730 ;
        RECT  7.265 2.310 8.700 2.730 ;
        RECT  7.095 2.265 7.265 2.730 ;
        RECT  5.750 2.310 7.095 2.730 ;
        RECT  5.580 2.265 5.750 2.730 ;
        RECT  4.390 2.310 5.580 2.730 ;
        RECT  4.220 2.265 4.390 2.730 ;
        RECT  3.790 2.310 4.220 2.730 ;
        RECT  3.620 2.215 3.790 2.730 ;
        RECT  3.095 2.310 3.620 2.730 ;
        RECT  2.925 2.215 3.095 2.730 ;
        RECT  1.575 2.310 2.925 2.730 ;
        RECT  1.405 2.265 1.575 2.730 ;
        RECT  0.605 2.310 1.405 2.730 ;
        RECT  0.435 2.185 0.605 2.730 ;
        RECT  0.000 2.310 0.435 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 12.040 2.520 ;
        LAYER M1 ;
        RECT  11.400 1.000 11.660 1.260 ;
        RECT  11.280 0.430 11.400 1.260 ;
        RECT  9.955 0.430 11.280 0.550 ;
        RECT  10.990 0.735 11.160 1.545 ;
        RECT  10.870 1.065 10.990 1.235 ;
        RECT  10.630 0.810 10.750 2.140 ;
        RECT  10.230 0.810 10.630 0.930 ;
        RECT  10.195 2.020 10.630 2.140 ;
        RECT  10.340 1.500 10.510 1.670 ;
        RECT  9.905 1.500 10.340 1.620 ;
        RECT  10.060 0.690 10.230 0.930 ;
        RECT  9.345 1.740 10.195 1.860 ;
        RECT  9.935 2.020 10.195 2.180 ;
        RECT  9.905 0.365 9.955 0.550 ;
        RECT  8.240 2.020 9.935 2.140 ;
        RECT  9.785 0.365 9.905 1.620 ;
        RECT  9.575 1.500 9.785 1.620 ;
        RECT  9.535 0.420 9.655 1.165 ;
        RECT  8.485 0.420 9.535 0.540 ;
        RECT  9.485 0.995 9.535 1.165 ;
        RECT  9.345 0.675 9.395 0.845 ;
        RECT  9.225 0.675 9.345 1.860 ;
        RECT  8.990 1.395 9.225 1.860 ;
        RECT  8.655 1.055 9.040 1.225 ;
        RECT  8.655 1.740 8.990 1.860 ;
        RECT  8.535 0.730 8.655 1.500 ;
        RECT  8.395 1.740 8.655 1.900 ;
        RECT  8.275 0.730 8.535 0.850 ;
        RECT  7.965 1.380 8.535 1.500 ;
        RECT  8.370 0.330 8.485 0.540 ;
        RECT  8.155 1.080 8.415 1.235 ;
        RECT  8.225 0.330 8.370 0.500 ;
        RECT  8.015 0.620 8.275 0.850 ;
        RECT  8.120 1.705 8.240 2.140 ;
        RECT  7.740 0.380 8.225 0.500 ;
        RECT  7.730 1.080 8.155 1.200 ;
        RECT  7.595 1.705 8.120 1.825 ;
        RECT  7.830 1.970 8.000 2.140 ;
        RECT  7.795 1.380 7.965 1.585 ;
        RECT  5.140 2.020 7.830 2.140 ;
        RECT  7.620 0.380 7.740 0.655 ;
        RECT  7.595 0.835 7.730 1.200 ;
        RECT  7.065 0.535 7.620 0.655 ;
        RECT  7.560 0.835 7.595 1.900 ;
        RECT  7.475 1.080 7.560 1.900 ;
        RECT  6.050 1.780 7.475 1.900 ;
        RECT  7.065 1.030 7.355 1.290 ;
        RECT  6.945 0.440 7.065 1.595 ;
        RECT  6.410 1.475 6.945 1.595 ;
        RECT  6.750 0.790 6.815 1.050 ;
        RECT  6.630 0.545 6.750 1.290 ;
        RECT  6.580 0.545 6.630 0.715 ;
        RECT  6.290 1.170 6.630 1.290 ;
        RECT  6.170 1.170 6.290 1.460 ;
        RECT  6.050 0.580 6.125 0.700 ;
        RECT  5.930 0.580 6.050 1.900 ;
        RECT  5.865 0.580 5.930 0.700 ;
        RECT  5.415 0.445 5.440 0.615 ;
        RECT  5.415 1.505 5.440 1.675 ;
        RECT  5.295 0.445 5.415 1.675 ;
        RECT  5.270 0.445 5.295 0.615 ;
        RECT  5.270 1.505 5.295 1.675 ;
        RECT  5.020 0.425 5.140 2.140 ;
        RECT  4.875 0.425 5.020 0.595 ;
        RECT  4.900 1.375 5.020 1.545 ;
        RECT  4.030 2.020 5.020 2.140 ;
        RECT  4.755 1.055 4.890 1.225 ;
        RECT  4.755 1.710 4.790 1.880 ;
        RECT  4.635 0.575 4.755 1.880 ;
        RECT  4.555 0.575 4.635 0.835 ;
        RECT  4.605 1.710 4.635 1.880 ;
        RECT  4.435 1.020 4.515 1.280 ;
        RECT  4.315 0.645 4.435 1.665 ;
        RECT  3.795 0.645 4.315 0.765 ;
        RECT  4.155 1.495 4.315 1.665 ;
        RECT  3.910 1.670 4.030 2.140 ;
        RECT  2.420 1.670 3.910 1.790 ;
        RECT  2.660 1.910 3.515 2.030 ;
        RECT  2.965 1.405 3.455 1.525 ;
        RECT  2.965 0.620 3.045 0.790 ;
        RECT  2.835 0.620 2.965 1.525 ;
        RECT  2.665 0.935 2.835 1.110 ;
        RECT  2.495 1.380 2.715 1.550 ;
        RECT  2.540 1.910 2.660 2.140 ;
        RECT  0.895 2.020 2.540 2.140 ;
        RECT  2.495 0.690 2.520 0.950 ;
        RECT  2.375 0.660 2.495 1.550 ;
        RECT  2.270 1.670 2.420 1.900 ;
        RECT  1.900 0.660 2.375 0.780 ;
        RECT  1.250 1.780 2.270 1.900 ;
        RECT  1.720 1.540 2.030 1.660 ;
        RECT  1.810 0.620 1.900 0.780 ;
        RECT  1.430 0.620 1.810 0.740 ;
        RECT  1.600 0.860 1.720 1.660 ;
        RECT  1.550 0.860 1.600 1.030 ;
        RECT  1.310 0.620 1.430 1.390 ;
        RECT  1.190 1.600 1.250 1.900 ;
        RECT  1.070 0.690 1.190 1.900 ;
        RECT  0.775 1.730 0.895 2.140 ;
        RECT  0.255 1.730 0.775 1.875 ;
        RECT  0.190 0.735 0.255 0.905 ;
        RECT  0.190 1.705 0.255 1.875 ;
        RECT  0.070 0.735 0.190 1.875 ;
    END
END SMDFFHQX2AD
MACRO SMDFFHQX4AD
    CLASS CORE ;
    FOREIGN SMDFFHQX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.115 0.770 1.375 ;
        END
        AntennaGateArea 0.072 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.365 0.905 3.765 1.025 ;
        RECT  3.245 0.590 3.365 1.025 ;
        RECT  3.110 0.590 3.245 0.710 ;
        RECT  2.990 0.380 3.110 0.710 ;
        RECT  1.100 0.380 2.990 0.500 ;
        RECT  0.960 0.350 1.100 0.500 ;
        RECT  0.840 0.350 0.960 0.560 ;
        RECT  0.490 0.440 0.840 0.560 ;
        RECT  0.350 0.440 0.490 0.815 ;
        RECT  0.160 0.440 0.350 0.560 ;
        END
        AntennaGateArea 0.138 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.915 0.780 4.035 1.330 ;
        RECT  3.665 1.160 3.915 1.330 ;
        RECT  3.075 1.160 3.665 1.280 ;
        RECT  2.955 1.020 3.075 1.280 ;
        END
        AntennaGateArea 0.1 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.555 1.005 13.650 1.515 ;
        RECT  13.385 0.400 13.555 2.145 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.635 1.100 1.890 1.375 ;
        END
        AntennaGateArea 0.143 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.300 0.865 5.545 1.200 ;
        END
        AntennaGateArea 0.143 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  5.905 0.910 6.275 1.120 ;
        END
        AntennaGateArea 0.191 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.915 -0.210 14.000 0.210 ;
        RECT  13.745 -0.210 13.915 0.795 ;
        RECT  13.005 -0.210 13.745 0.210 ;
        RECT  12.835 -0.210 13.005 0.255 ;
        RECT  11.035 -0.210 12.835 0.210 ;
        RECT  10.865 -0.210 11.035 0.255 ;
        RECT  10.275 -0.210 10.865 0.210 ;
        RECT  10.105 -0.210 10.275 0.255 ;
        RECT  9.305 -0.210 10.105 0.210 ;
        RECT  9.135 -0.210 9.305 0.255 ;
        RECT  7.960 -0.210 9.135 0.210 ;
        RECT  7.790 -0.210 7.960 0.255 ;
        RECT  6.720 -0.210 7.790 0.210 ;
        RECT  6.550 -0.210 6.720 0.255 ;
        RECT  5.685 -0.210 6.550 0.210 ;
        RECT  5.515 -0.210 5.685 0.255 ;
        RECT  4.215 -0.210 5.515 0.210 ;
        RECT  4.045 -0.210 4.215 0.255 ;
        RECT  3.455 -0.210 4.045 0.210 ;
        RECT  3.285 -0.210 3.455 0.255 ;
        RECT  2.130 -0.210 3.285 0.210 ;
        RECT  1.960 -0.210 2.130 0.255 ;
        RECT  0.590 -0.210 1.960 0.210 ;
        RECT  0.420 -0.210 0.590 0.320 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  13.905 2.310 14.000 2.730 ;
        RECT  13.770 1.400 13.905 2.730 ;
        RECT  13.195 2.310 13.770 2.730 ;
        RECT  13.025 1.835 13.195 2.730 ;
        RECT  12.635 2.310 13.025 2.730 ;
        RECT  12.465 1.730 12.635 2.730 ;
        RECT  10.985 2.310 12.465 2.730 ;
        RECT  10.815 2.265 10.985 2.730 ;
        RECT  10.215 2.310 10.815 2.730 ;
        RECT  10.045 2.265 10.215 2.730 ;
        RECT  9.285 2.310 10.045 2.730 ;
        RECT  9.115 2.265 9.285 2.730 ;
        RECT  8.005 2.310 9.115 2.730 ;
        RECT  7.835 2.265 8.005 2.730 ;
        RECT  7.210 2.310 7.835 2.730 ;
        RECT  7.040 2.265 7.210 2.730 ;
        RECT  6.240 2.310 7.040 2.730 ;
        RECT  6.070 2.265 6.240 2.730 ;
        RECT  5.685 2.310 6.070 2.730 ;
        RECT  5.515 2.265 5.685 2.730 ;
        RECT  4.215 2.310 5.515 2.730 ;
        RECT  4.045 2.265 4.215 2.730 ;
        RECT  3.670 2.310 4.045 2.730 ;
        RECT  3.500 2.265 3.670 2.730 ;
        RECT  2.910 2.310 3.500 2.730 ;
        RECT  2.740 2.265 2.910 2.730 ;
        RECT  1.560 2.310 2.740 2.730 ;
        RECT  1.390 2.265 1.560 2.730 ;
        RECT  0.590 2.310 1.390 2.730 ;
        RECT  0.420 2.085 0.590 2.730 ;
        RECT  0.000 2.310 0.420 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 14.000 2.520 ;
        LAYER M1 ;
        RECT  13.155 1.050 13.205 1.220 ;
        RECT  13.035 0.380 13.155 1.220 ;
        RECT  12.240 0.380 13.035 0.500 ;
        RECT  12.715 0.735 12.885 1.545 ;
        RECT  12.400 1.115 12.715 1.285 ;
        RECT  12.280 0.620 12.375 0.790 ;
        RECT  12.160 0.620 12.280 2.140 ;
        RECT  12.040 0.330 12.240 0.500 ;
        RECT  12.005 1.965 12.160 2.140 ;
        RECT  11.980 0.330 12.040 1.605 ;
        RECT  9.665 2.020 12.005 2.140 ;
        RECT  11.920 0.380 11.980 1.605 ;
        RECT  11.395 0.380 11.920 0.500 ;
        RECT  11.805 1.435 11.920 1.605 ;
        RECT  11.255 1.485 11.805 1.605 ;
        RECT  11.660 0.630 11.800 0.750 ;
        RECT  11.540 0.630 11.660 1.325 ;
        RECT  11.445 1.730 11.615 1.900 ;
        RECT  10.685 1.205 11.540 1.325 ;
        RECT  10.685 1.780 11.445 1.900 ;
        RECT  11.275 0.380 11.395 0.720 ;
        RECT  11.225 0.550 11.275 0.720 ;
        RECT  11.085 1.485 11.255 1.655 ;
        RECT  10.935 0.960 11.180 1.080 ;
        RECT  10.815 0.380 10.935 1.080 ;
        RECT  7.805 0.380 10.815 0.500 ;
        RECT  10.680 1.205 10.685 1.900 ;
        RECT  10.560 0.635 10.680 1.900 ;
        RECT  10.485 0.635 10.560 0.805 ;
        RECT  10.435 1.470 10.560 1.900 ;
        RECT  9.800 1.780 10.435 1.900 ;
        RECT  10.135 0.975 10.430 1.145 ;
        RECT  10.015 0.740 10.135 1.545 ;
        RECT  9.690 0.740 10.015 0.860 ;
        RECT  8.645 1.425 10.015 1.545 ;
        RECT  9.430 0.660 9.690 0.860 ;
        RECT  9.545 1.740 9.665 2.140 ;
        RECT  8.355 1.740 9.545 1.860 ;
        RECT  8.355 1.110 9.490 1.230 ;
        RECT  8.655 0.740 9.430 0.860 ;
        RECT  8.300 1.980 8.820 2.190 ;
        RECT  8.485 0.620 8.655 0.860 ;
        RECT  8.475 1.375 8.645 1.545 ;
        RECT  8.235 0.850 8.355 1.860 ;
        RECT  4.920 1.980 8.300 2.100 ;
        RECT  8.190 0.850 8.235 0.970 ;
        RECT  6.515 1.740 8.235 1.860 ;
        RECT  7.930 0.820 8.190 0.970 ;
        RECT  7.805 1.125 8.115 1.265 ;
        RECT  7.685 0.380 7.805 1.580 ;
        RECT  7.370 0.380 7.685 0.550 ;
        RECT  6.905 1.460 7.685 1.580 ;
        RECT  7.100 0.850 7.480 1.130 ;
        RECT  7.050 0.380 7.100 1.130 ;
        RECT  6.930 0.380 7.050 0.970 ;
        RECT  5.785 0.380 6.930 0.500 ;
        RECT  6.785 1.140 6.905 1.580 ;
        RECT  6.645 1.140 6.785 1.260 ;
        RECT  6.395 0.620 6.515 1.860 ;
        RECT  6.125 0.620 6.395 0.740 ;
        RECT  5.785 1.450 5.990 1.620 ;
        RECT  5.665 0.380 5.785 1.620 ;
        RECT  5.165 0.470 5.305 0.640 ;
        RECT  5.165 1.380 5.305 1.810 ;
        RECT  5.135 0.470 5.165 1.810 ;
        RECT  5.045 0.470 5.135 1.500 ;
        RECT  4.780 0.360 4.920 2.100 ;
        RECT  3.805 1.980 4.780 2.100 ;
        RECT  4.540 0.515 4.660 1.860 ;
        RECT  4.425 0.515 4.540 0.685 ;
        RECT  4.400 1.740 4.540 1.860 ;
        RECT  4.305 0.990 4.360 1.250 ;
        RECT  4.210 0.540 4.305 1.615 ;
        RECT  4.185 0.540 4.210 1.665 ;
        RECT  3.630 0.540 4.185 0.660 ;
        RECT  4.040 1.495 4.185 1.665 ;
        RECT  3.685 1.660 3.805 2.100 ;
        RECT  3.005 1.660 3.685 1.780 ;
        RECT  3.240 1.920 3.410 2.140 ;
        RECT  2.835 1.420 3.335 1.540 ;
        RECT  1.145 2.020 3.240 2.140 ;
        RECT  2.885 1.660 3.005 1.900 ;
        RECT  1.195 1.780 2.885 1.900 ;
        RECT  2.715 0.660 2.835 1.540 ;
        RECT  2.650 0.660 2.715 0.830 ;
        RECT  2.570 1.065 2.715 1.235 ;
        RECT  2.475 1.380 2.595 1.640 ;
        RECT  2.435 1.380 2.475 1.500 ;
        RECT  2.315 0.620 2.435 1.500 ;
        RECT  1.390 0.620 2.315 0.740 ;
        RECT  2.025 0.860 2.145 1.660 ;
        RECT  1.510 0.860 2.025 0.980 ;
        RECT  1.775 1.540 2.025 1.660 ;
        RECT  1.270 0.620 1.390 1.395 ;
        RECT  1.150 1.550 1.195 1.900 ;
        RECT  1.030 0.680 1.150 1.900 ;
        RECT  0.910 2.020 1.145 2.170 ;
        RECT  0.885 1.735 0.910 2.170 ;
        RECT  0.790 1.735 0.885 2.140 ;
        RECT  0.255 1.735 0.790 1.855 ;
        RECT  0.205 1.585 0.255 1.855 ;
        RECT  0.205 0.680 0.230 0.940 ;
        RECT  0.085 0.680 0.205 1.855 ;
    END
END SMDFFHQX4AD
MACRO SMDFFHQX8AD
    CLASS CORE ;
    FOREIGN SMDFFHQX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.440 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.690 1.115 0.770 1.375 ;
        RECT  0.570 1.010 0.690 1.375 ;
        RECT  0.350 1.115 0.570 1.375 ;
        END
        AntennaGateArea 0.136 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.970 0.905 5.315 1.025 ;
        RECT  4.830 0.380 4.970 1.025 ;
        RECT  0.375 0.380 4.830 0.500 ;
        RECT  0.205 0.380 0.375 0.550 ;
        END
        AntennaGateArea 0.165 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.465 0.780 5.585 1.330 ;
        RECT  5.065 1.160 5.465 1.330 ;
        RECT  4.665 1.160 5.065 1.280 ;
        RECT  4.545 1.020 4.665 1.280 ;
        END
        AntennaGateArea 0.12 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  19.825 0.400 19.995 2.145 ;
        RECT  19.275 1.005 19.825 1.515 ;
        RECT  19.105 0.400 19.275 2.145 ;
        END
        AntennaDiffArea 0.844 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.705 0.910 2.285 1.085 ;
        END
        AntennaGateArea 0.274 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.585 0.910 8.095 1.145 ;
        END
        AntennaGateArea 0.274 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  9.740 0.905 10.335 1.075 ;
        END
        AntennaGateArea 0.344 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  20.355 -0.210 20.440 0.210 ;
        RECT  20.185 -0.210 20.355 0.795 ;
        RECT  19.635 -0.210 20.185 0.210 ;
        RECT  19.465 -0.210 19.635 0.795 ;
        RECT  18.715 -0.210 19.465 0.210 ;
        RECT  18.545 -0.210 18.715 0.255 ;
        RECT  15.995 -0.210 18.545 0.210 ;
        RECT  15.825 -0.210 15.995 0.255 ;
        RECT  15.235 -0.210 15.825 0.210 ;
        RECT  15.065 -0.210 15.235 0.255 ;
        RECT  14.475 -0.210 15.065 0.210 ;
        RECT  14.305 -0.210 14.475 0.255 ;
        RECT  13.570 -0.210 14.305 0.210 ;
        RECT  13.400 -0.210 13.570 0.255 ;
        RECT  12.285 -0.210 13.400 0.210 ;
        RECT  12.025 -0.210 12.285 0.380 ;
        RECT  11.150 -0.210 12.025 0.210 ;
        RECT  10.980 -0.210 11.150 0.255 ;
        RECT  10.375 -0.210 10.980 0.210 ;
        RECT  10.205 -0.210 10.375 0.255 ;
        RECT  9.615 -0.210 10.205 0.210 ;
        RECT  9.445 -0.210 9.615 0.255 ;
        RECT  9.275 -0.210 9.445 0.210 ;
        RECT  9.105 -0.210 9.275 0.255 ;
        RECT  8.330 -0.210 9.105 0.210 ;
        RECT  8.160 -0.210 8.330 0.760 ;
        RECT  7.610 -0.210 8.160 0.210 ;
        RECT  7.440 -0.210 7.610 0.450 ;
        RECT  5.840 -0.210 7.440 0.210 ;
        RECT  5.670 -0.210 5.840 0.255 ;
        RECT  5.170 -0.210 5.670 0.210 ;
        RECT  5.000 -0.210 5.170 0.255 ;
        RECT  3.890 -0.210 5.000 0.210 ;
        RECT  3.720 -0.210 3.890 0.255 ;
        RECT  2.500 -0.210 3.720 0.210 ;
        RECT  2.330 -0.210 2.500 0.255 ;
        RECT  1.735 -0.210 2.330 0.210 ;
        RECT  1.565 -0.210 1.735 0.255 ;
        RECT  0.590 -0.210 1.565 0.210 ;
        RECT  0.420 -0.210 0.590 0.255 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  20.355 2.310 20.440 2.730 ;
        RECT  20.185 1.445 20.355 2.730 ;
        RECT  19.635 2.310 20.185 2.730 ;
        RECT  19.465 1.785 19.635 2.730 ;
        RECT  18.915 2.310 19.465 2.730 ;
        RECT  18.745 1.835 18.915 2.730 ;
        RECT  18.340 2.310 18.745 2.730 ;
        RECT  18.170 1.725 18.340 2.730 ;
        RECT  15.995 2.310 18.170 2.730 ;
        RECT  15.825 2.265 15.995 2.730 ;
        RECT  15.235 2.310 15.825 2.730 ;
        RECT  15.065 2.265 15.235 2.730 ;
        RECT  14.475 2.310 15.065 2.730 ;
        RECT  14.305 2.265 14.475 2.730 ;
        RECT  13.520 2.310 14.305 2.730 ;
        RECT  13.350 1.930 13.520 2.730 ;
        RECT  12.285 2.310 13.350 2.730 ;
        RECT  12.025 2.130 12.285 2.730 ;
        RECT  11.385 2.310 12.025 2.730 ;
        RECT  11.125 2.130 11.385 2.730 ;
        RECT  10.030 2.310 11.125 2.730 ;
        RECT  9.860 2.265 10.030 2.730 ;
        RECT  9.000 2.310 9.860 2.730 ;
        RECT  8.830 2.265 9.000 2.730 ;
        RECT  8.240 2.310 8.830 2.730 ;
        RECT  8.070 2.265 8.240 2.730 ;
        RECT  7.480 2.310 8.070 2.730 ;
        RECT  7.310 2.265 7.480 2.730 ;
        RECT  5.220 2.310 7.310 2.730 ;
        RECT  5.050 2.265 5.220 2.730 ;
        RECT  4.460 2.310 5.050 2.730 ;
        RECT  4.290 2.265 4.460 2.730 ;
        RECT  2.500 2.310 4.290 2.730 ;
        RECT  2.330 2.265 2.500 2.730 ;
        RECT  1.740 2.310 2.330 2.730 ;
        RECT  1.570 2.265 1.740 2.730 ;
        RECT  0.590 2.310 1.570 2.730 ;
        RECT  0.420 1.965 0.590 2.730 ;
        RECT  0.000 2.310 0.420 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 20.440 2.520 ;
        LAYER M1 ;
        RECT  18.875 1.050 18.925 1.220 ;
        RECT  18.755 0.380 18.875 1.220 ;
        RECT  17.895 0.380 18.755 0.500 ;
        RECT  18.435 0.735 18.605 1.545 ;
        RECT  18.125 1.115 18.435 1.285 ;
        RECT  17.965 0.630 18.135 0.750 ;
        RECT  17.845 0.630 17.965 2.190 ;
        RECT  17.710 0.330 17.895 0.500 ;
        RECT  17.705 2.020 17.845 2.190 ;
        RECT  17.635 0.330 17.710 1.715 ;
        RECT  13.945 2.020 17.705 2.140 ;
        RECT  17.590 0.380 17.635 1.715 ;
        RECT  16.150 0.380 17.590 0.500 ;
        RECT  17.540 1.485 17.590 1.715 ;
        RECT  16.265 1.485 17.540 1.605 ;
        RECT  17.300 0.620 17.470 0.790 ;
        RECT  17.175 1.730 17.345 1.900 ;
        RECT  16.675 0.620 17.300 0.740 ;
        RECT  15.615 1.780 17.175 1.900 ;
        RECT  16.555 0.620 16.675 1.365 ;
        RECT  16.010 0.620 16.555 0.740 ;
        RECT  15.615 1.245 16.555 1.365 ;
        RECT  16.095 1.485 16.265 1.655 ;
        RECT  15.975 0.935 16.145 1.105 ;
        RECT  15.890 0.425 16.010 0.740 ;
        RECT  15.760 0.935 15.975 1.055 ;
        RECT  14.855 0.425 15.890 0.545 ;
        RECT  15.640 0.735 15.760 1.055 ;
        RECT  14.565 0.735 15.640 0.855 ;
        RECT  15.495 1.245 15.615 1.900 ;
        RECT  15.445 1.470 15.495 1.900 ;
        RECT  14.855 1.780 15.445 1.900 ;
        RECT  14.325 0.975 15.325 1.145 ;
        RECT  14.685 0.375 14.855 0.545 ;
        RECT  14.685 1.470 14.855 1.900 ;
        RECT  14.090 1.780 14.685 1.900 ;
        RECT  14.445 0.380 14.565 0.855 ;
        RECT  14.100 0.380 14.445 0.500 ;
        RECT  14.205 0.750 14.325 1.470 ;
        RECT  13.980 0.750 14.205 0.870 ;
        RECT  12.880 1.350 14.205 1.470 ;
        RECT  13.840 0.355 14.100 0.500 ;
        RECT  13.720 0.645 13.980 0.870 ;
        RECT  13.775 1.640 13.945 2.140 ;
        RECT  12.545 0.380 13.840 0.500 ;
        RECT  10.660 1.640 13.775 1.760 ;
        RECT  12.925 0.750 13.720 0.870 ;
        RECT  12.655 2.070 13.055 2.190 ;
        RECT  12.665 0.630 12.925 0.870 ;
        RECT  12.710 1.350 12.880 1.520 ;
        RECT  11.610 1.350 12.710 1.470 ;
        RECT  11.655 0.750 12.665 0.870 ;
        RECT  12.535 1.890 12.655 2.190 ;
        RECT  12.425 0.380 12.545 0.620 ;
        RECT  11.775 1.890 12.535 2.010 ;
        RECT  11.895 0.500 12.425 0.620 ;
        RECT  11.775 0.380 11.895 0.620 ;
        RECT  9.210 0.380 11.775 0.500 ;
        RECT  11.515 1.890 11.775 2.190 ;
        RECT  11.395 0.630 11.655 0.870 ;
        RECT  11.440 1.350 11.610 1.520 ;
        RECT  10.835 1.890 11.515 2.010 ;
        RECT  10.660 0.990 11.440 1.160 ;
        RECT  10.715 1.890 10.835 2.140 ;
        RECT  10.660 0.620 10.815 0.740 ;
        RECT  9.325 2.020 10.715 2.140 ;
        RECT  10.540 0.620 10.660 1.760 ;
        RECT  10.490 1.330 10.540 1.760 ;
        RECT  9.620 0.620 10.040 0.740 ;
        RECT  9.620 1.370 9.720 1.800 ;
        RECT  9.500 0.620 9.620 1.800 ;
        RECT  8.710 0.995 9.500 1.165 ;
        RECT  9.210 1.305 9.380 1.735 ;
        RECT  9.205 1.890 9.325 2.140 ;
        RECT  9.090 0.380 9.210 0.715 ;
        RECT  8.620 1.305 9.210 1.425 ;
        RECT  6.850 1.890 9.205 2.010 ;
        RECT  8.895 0.595 9.090 0.715 ;
        RECT  8.570 0.595 8.895 0.765 ;
        RECT  8.570 1.305 8.620 1.735 ;
        RECT  8.450 0.595 8.570 1.735 ;
        RECT  7.800 0.470 7.970 0.700 ;
        RECT  7.690 1.330 7.860 1.760 ;
        RECT  7.455 0.580 7.800 0.700 ;
        RECT  7.455 1.640 7.690 1.760 ;
        RECT  7.335 0.580 7.455 1.760 ;
        RECT  6.490 1.640 7.335 1.760 ;
        RECT  7.140 0.650 7.190 0.820 ;
        RECT  7.140 1.345 7.190 1.515 ;
        RECT  7.020 0.650 7.140 1.515 ;
        RECT  6.775 1.020 7.020 1.280 ;
        RECT  6.680 0.380 6.850 0.640 ;
        RECT  6.680 1.890 6.850 2.060 ;
        RECT  6.130 0.380 6.680 0.500 ;
        RECT  6.130 1.890 6.680 2.010 ;
        RECT  6.370 0.640 6.490 1.760 ;
        RECT  6.320 0.640 6.370 0.810 ;
        RECT  6.320 1.410 6.370 1.580 ;
        RECT  6.010 0.380 6.130 2.010 ;
        RECT  5.960 0.610 6.010 0.780 ;
        RECT  5.960 1.380 6.010 2.010 ;
        RECT  5.355 1.890 5.960 2.010 ;
        RECT  5.840 0.900 5.890 1.160 ;
        RECT  5.790 0.540 5.840 1.615 ;
        RECT  5.720 0.540 5.790 1.665 ;
        RECT  5.245 0.540 5.720 0.660 ;
        RECT  5.620 1.495 5.720 1.665 ;
        RECT  5.235 1.660 5.355 2.010 ;
        RECT  4.555 1.660 5.235 1.780 ;
        RECT  4.790 1.920 4.960 2.140 ;
        RECT  4.425 1.420 4.885 1.540 ;
        RECT  0.835 2.020 4.790 2.140 ;
        RECT  4.435 1.660 4.555 1.900 ;
        RECT  4.425 0.660 4.520 0.830 ;
        RECT  3.215 1.780 4.435 1.900 ;
        RECT  4.305 0.660 4.425 1.540 ;
        RECT  4.150 1.045 4.305 1.215 ;
        RECT  4.015 0.660 4.180 0.830 ;
        RECT  4.015 1.380 4.055 1.640 ;
        RECT  3.895 0.660 4.015 1.640 ;
        RECT  3.645 1.210 3.895 1.380 ;
        RECT  3.510 1.485 3.560 1.655 ;
        RECT  3.510 0.620 3.550 0.805 ;
        RECT  3.390 0.620 3.510 1.655 ;
        RECT  3.380 0.620 3.390 0.805 ;
        RECT  2.790 0.620 3.380 0.740 ;
        RECT  3.095 0.860 3.215 1.900 ;
        RECT  2.955 0.860 3.095 0.980 ;
        RECT  3.030 1.730 3.095 1.900 ;
        RECT  1.220 1.780 3.030 1.900 ;
        RECT  2.790 1.400 2.840 1.655 ;
        RECT  2.670 0.620 2.790 1.655 ;
        RECT  2.620 0.620 2.670 0.805 ;
        RECT  2.120 1.400 2.670 1.520 ;
        RECT  1.900 0.620 2.620 0.740 ;
        RECT  1.950 1.400 2.120 1.570 ;
        RECT  1.145 0.715 1.240 0.885 ;
        RECT  1.145 1.470 1.220 1.900 ;
        RECT  1.070 0.715 1.145 1.900 ;
        RECT  1.025 0.750 1.070 1.900 ;
        RECT  0.715 1.675 0.835 2.140 ;
        RECT  0.255 1.675 0.715 1.795 ;
        RECT  0.205 0.715 0.255 0.885 ;
        RECT  0.205 1.455 0.255 1.795 ;
        RECT  0.085 0.715 0.205 1.795 ;
    END
END SMDFFHQX8AD
MACRO TBUFX12AD
    CLASS CORE ;
    FOREIGN TBUFX12AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  5.500 0.340 5.670 0.770 ;
        RECT  5.310 0.570 5.500 0.770 ;
        RECT  5.120 0.570 5.310 2.160 ;
        RECT  4.950 0.570 5.120 1.675 ;
        RECT  4.780 0.340 4.950 1.675 ;
        RECT  4.585 0.570 4.780 1.675 ;
        RECT  4.495 0.570 4.585 1.970 ;
        RECT  4.230 0.570 4.495 0.710 ;
        RECT  4.415 1.500 4.495 1.970 ;
        RECT  3.880 1.500 4.415 1.675 ;
        RECT  4.060 0.340 4.230 0.770 ;
        RECT  3.505 0.570 4.060 0.710 ;
        RECT  3.680 1.500 3.880 2.160 ;
        RECT  3.335 0.340 3.505 0.770 ;
        END
        AntennaDiffArea 1.198 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.425 0.430 1.545 ;
        RECT  0.070 1.425 0.210 1.655 ;
        END
        AntennaGateArea 0.2074 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.100 1.145 2.895 1.375 ;
        END
        AntennaGateArea 0.372 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.355 -0.210 5.880 0.210 ;
        RECT  5.095 -0.210 5.355 0.430 ;
        RECT  4.635 -0.210 5.095 0.210 ;
        RECT  4.375 -0.210 4.635 0.430 ;
        RECT  3.915 -0.210 4.375 0.210 ;
        RECT  3.645 -0.210 3.915 0.430 ;
        RECT  3.155 -0.210 3.645 0.210 ;
        RECT  2.895 -0.210 3.155 0.640 ;
        RECT  2.435 -0.210 2.895 0.210 ;
        RECT  2.175 -0.210 2.435 0.640 ;
        RECT  0.865 -0.210 2.175 0.210 ;
        RECT  0.480 -0.210 0.865 0.760 ;
        RECT  0.000 -0.210 0.480 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.665 2.310 5.880 2.730 ;
        RECT  5.495 1.520 5.665 2.730 ;
        RECT  4.945 2.310 5.495 2.730 ;
        RECT  4.775 1.845 4.945 2.730 ;
        RECT  4.225 2.310 4.775 2.730 ;
        RECT  4.055 1.845 4.225 2.730 ;
        RECT  3.510 2.310 4.055 2.730 ;
        RECT  3.340 1.640 3.510 2.730 ;
        RECT  2.805 2.310 3.340 2.730 ;
        RECT  2.635 1.800 2.805 2.730 ;
        RECT  2.085 2.310 2.635 2.730 ;
        RECT  1.910 1.845 2.085 2.730 ;
        RECT  0.265 2.310 1.910 2.730 ;
        RECT  0.095 1.795 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.880 2.520 ;
        LAYER M1 ;
        RECT  3.240 0.905 4.370 1.025 ;
        RECT  3.180 1.210 4.330 1.330 ;
        RECT  3.115 0.855 3.240 1.025 ;
        RECT  3.020 1.210 3.180 2.160 ;
        RECT  2.750 0.855 3.115 0.975 ;
        RECT  2.475 1.545 3.020 1.680 ;
        RECT  2.580 0.400 2.750 0.975 ;
        RECT  2.045 0.855 2.580 0.975 ;
        RECT  2.245 1.545 2.475 2.050 ;
        RECT  1.725 1.545 2.245 1.680 ;
        RECT  1.845 0.435 2.045 0.975 ;
        RECT  1.255 0.435 1.845 0.575 ;
        RECT  1.670 1.545 1.725 2.110 ;
        RECT  1.500 0.775 1.670 2.110 ;
        RECT  0.985 1.990 1.500 2.110 ;
        RECT  1.255 0.785 1.375 1.825 ;
        RECT  1.240 0.435 1.255 1.825 ;
        RECT  1.085 0.435 1.240 1.060 ;
        RECT  1.175 1.655 1.240 1.825 ;
        RECT  0.670 1.290 1.105 1.485 ;
        RECT  0.815 1.665 0.985 2.110 ;
        RECT  0.550 1.185 0.670 2.055 ;
        RECT  0.240 1.185 0.550 1.305 ;
        RECT  0.465 1.885 0.550 2.055 ;
        RECT  0.120 0.460 0.240 1.305 ;
    END
END TBUFX12AD
MACRO TBUFX16AD
    CLASS CORE ;
    FOREIGN TBUFX16AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  6.240 0.345 6.410 0.775 ;
        RECT  6.110 0.570 6.240 0.775 ;
        RECT  6.045 0.570 6.110 1.675 ;
        RECT  5.875 0.570 6.045 1.930 ;
        RECT  5.690 0.570 5.875 1.675 ;
        RECT  5.520 0.340 5.690 1.675 ;
        RECT  5.370 0.570 5.520 1.675 ;
        RECT  4.970 0.570 5.370 0.710 ;
        RECT  5.330 1.500 5.370 1.675 ;
        RECT  5.140 1.500 5.330 2.160 ;
        RECT  4.605 1.500 5.140 1.675 ;
        RECT  4.800 0.340 4.970 0.770 ;
        RECT  3.530 0.570 4.800 0.710 ;
        RECT  4.435 1.500 4.605 1.970 ;
        RECT  3.900 1.500 4.435 1.675 ;
        RECT  3.700 1.500 3.900 2.160 ;
        RECT  3.360 0.340 3.530 0.770 ;
        END
        AntennaDiffArea 1.585 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.425 0.430 1.545 ;
        RECT  0.070 1.425 0.210 1.655 ;
        END
        AntennaGateArea 0.268 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.510 1.235 3.230 1.375 ;
        RECT  2.190 1.145 2.510 1.375 ;
        END
        AntennaGateArea 0.475 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.095 -0.210 6.720 0.210 ;
        RECT  5.835 -0.210 6.095 0.430 ;
        RECT  5.375 -0.210 5.835 0.210 ;
        RECT  5.115 -0.210 5.375 0.430 ;
        RECT  4.655 -0.210 5.115 0.210 ;
        RECT  4.395 -0.210 4.655 0.430 ;
        RECT  3.935 -0.210 4.395 0.210 ;
        RECT  3.675 -0.210 3.935 0.430 ;
        RECT  3.210 -0.210 3.675 0.210 ;
        RECT  2.950 -0.210 3.210 0.665 ;
        RECT  2.490 -0.210 2.950 0.210 ;
        RECT  2.230 -0.210 2.490 0.690 ;
        RECT  0.900 -0.210 2.230 0.210 ;
        RECT  0.440 -0.210 0.900 0.880 ;
        RECT  0.000 -0.210 0.440 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.405 2.310 6.720 2.730 ;
        RECT  6.235 1.845 6.405 2.730 ;
        RECT  5.685 2.310 6.235 2.730 ;
        RECT  5.515 1.800 5.685 2.730 ;
        RECT  4.965 2.310 5.515 2.730 ;
        RECT  4.795 1.845 4.965 2.730 ;
        RECT  4.245 2.310 4.795 2.730 ;
        RECT  4.075 1.845 4.245 2.730 ;
        RECT  3.530 2.310 4.075 2.730 ;
        RECT  3.360 1.800 3.530 2.730 ;
        RECT  2.805 2.310 3.360 2.730 ;
        RECT  2.635 1.800 2.805 2.730 ;
        RECT  2.085 2.310 2.635 2.730 ;
        RECT  1.910 1.845 2.085 2.730 ;
        RECT  0.265 2.310 1.910 2.730 ;
        RECT  0.095 1.795 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.720 2.520 ;
        LAYER M1 ;
        RECT  3.570 1.210 5.240 1.330 ;
        RECT  3.320 0.905 5.080 1.050 ;
        RECT  3.435 1.210 3.570 1.680 ;
        RECT  3.180 1.545 3.435 1.680 ;
        RECT  2.805 0.905 3.320 1.025 ;
        RECT  2.980 1.545 3.180 2.160 ;
        RECT  2.475 1.545 2.980 1.680 ;
        RECT  2.635 0.435 2.805 1.025 ;
        RECT  2.085 0.905 2.635 1.025 ;
        RECT  2.245 1.545 2.475 2.050 ;
        RECT  1.725 1.545 2.245 1.680 ;
        RECT  1.915 0.405 2.085 1.025 ;
        RECT  1.400 0.405 1.915 0.525 ;
        RECT  1.555 0.695 1.725 2.110 ;
        RECT  0.985 1.975 1.555 2.110 ;
        RECT  1.265 0.405 1.400 1.825 ;
        RECT  1.175 0.405 1.265 0.865 ;
        RECT  1.175 1.655 1.265 1.825 ;
        RECT  0.670 1.245 1.070 1.505 ;
        RECT  0.815 1.665 0.985 2.110 ;
        RECT  0.550 1.185 0.670 2.055 ;
        RECT  0.240 1.185 0.550 1.305 ;
        RECT  0.465 1.885 0.550 2.055 ;
        RECT  0.120 0.530 0.240 1.305 ;
    END
END TBUFX16AD
MACRO TBUFX1AD
    CLASS CORE ;
    FOREIGN TBUFX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.280 0.355 2.450 2.115 ;
        RECT  2.215 0.355 2.280 0.525 ;
        END
        AntennaDiffArea 0.206 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.115 0.540 1.285 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.0888 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.620 1.145 1.890 1.375 ;
        END
        AntennaGateArea 0.0419 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.070 -0.210 2.520 0.210 ;
        RECT  1.810 -0.210 2.070 0.500 ;
        RECT  0.690 -0.210 1.810 0.210 ;
        RECT  0.570 -0.210 0.690 0.620 ;
        RECT  0.000 -0.210 0.570 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.080 2.310 2.520 2.730 ;
        RECT  1.820 1.740 2.080 2.730 ;
        RECT  0.245 2.310 1.820 2.730 ;
        RECT  0.095 1.670 0.245 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.110 0.710 2.150 0.970 ;
        RECT  2.030 1.255 2.150 1.620 ;
        RECT  1.990 0.640 2.110 0.970 ;
        RECT  1.630 1.500 2.030 1.620 ;
        RECT  1.690 0.640 1.990 0.760 ;
        RECT  1.570 0.380 1.690 0.760 ;
        RECT  1.500 0.880 1.680 1.000 ;
        RECT  1.510 1.500 1.630 2.130 ;
        RECT  1.430 0.380 1.570 0.550 ;
        RECT  1.500 1.500 1.510 1.620 ;
        RECT  0.420 2.010 1.510 2.130 ;
        RECT  1.380 0.880 1.500 1.620 ;
        RECT  1.250 0.430 1.430 0.550 ;
        RECT  1.250 1.720 1.285 1.890 ;
        RECT  1.130 0.430 1.250 1.890 ;
        RECT  0.860 0.430 1.130 0.550 ;
        RECT  1.095 1.720 1.130 1.890 ;
        RECT  0.900 1.500 0.965 1.670 ;
        RECT  0.780 0.750 0.900 1.670 ;
        RECT  0.450 0.750 0.780 0.875 ;
        RECT  0.490 1.410 0.780 1.670 ;
        RECT  0.330 0.430 0.450 0.875 ;
        RECT  0.130 0.430 0.330 0.550 ;
    END
END TBUFX1AD
MACRO TBUFX20AD
    CLASS CORE ;
    FOREIGN TBUFX20AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  7.865 0.570 8.070 1.675 ;
        RECT  7.860 0.570 7.865 1.930 ;
        RECT  7.695 0.345 7.860 1.930 ;
        RECT  7.690 0.345 7.695 1.675 ;
        RECT  7.295 0.570 7.690 1.675 ;
        RECT  7.140 0.570 7.295 0.710 ;
        RECT  7.145 1.500 7.295 1.675 ;
        RECT  6.975 1.500 7.145 1.930 ;
        RECT  6.970 0.345 7.140 0.775 ;
        RECT  6.430 1.500 6.975 1.675 ;
        RECT  6.420 0.570 6.970 0.710 ;
        RECT  6.240 1.500 6.430 2.160 ;
        RECT  6.250 0.345 6.420 0.775 ;
        RECT  5.700 0.570 6.250 0.710 ;
        RECT  5.705 1.500 6.240 1.675 ;
        RECT  5.535 1.500 5.705 1.970 ;
        RECT  5.530 0.345 5.700 0.775 ;
        RECT  5.000 1.500 5.535 1.675 ;
        RECT  4.980 0.570 5.530 0.710 ;
        RECT  4.800 1.500 5.000 2.160 ;
        RECT  4.810 0.345 4.980 0.775 ;
        RECT  4.255 0.570 4.810 0.710 ;
        RECT  4.085 0.345 4.255 0.775 ;
        END
        AntennaDiffArea 1.968 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.385 1.145 1.835 1.375 ;
        END
        AntennaGateArea 0.3348 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.065 1.220 3.965 1.375 ;
        RECT  2.820 1.145 3.065 1.375 ;
        END
        AntennaGateArea 0.5866 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.270 -0.210 8.400 0.210 ;
        RECT  8.010 -0.210 8.270 0.415 ;
        RECT  7.550 -0.210 8.010 0.210 ;
        RECT  7.280 -0.210 7.550 0.415 ;
        RECT  6.830 -0.210 7.280 0.210 ;
        RECT  6.560 -0.210 6.830 0.415 ;
        RECT  6.110 -0.210 6.560 0.210 ;
        RECT  5.840 -0.210 6.110 0.415 ;
        RECT  5.390 -0.210 5.840 0.210 ;
        RECT  5.120 -0.210 5.390 0.415 ;
        RECT  4.665 -0.210 5.120 0.210 ;
        RECT  4.405 -0.210 4.665 0.390 ;
        RECT  3.895 -0.210 4.405 0.210 ;
        RECT  3.725 -0.210 3.895 0.715 ;
        RECT  3.155 -0.210 3.725 0.210 ;
        RECT  2.985 -0.210 3.155 0.715 ;
        RECT  2.435 -0.210 2.985 0.210 ;
        RECT  2.265 -0.210 2.435 0.455 ;
        RECT  1.740 -0.210 2.265 0.210 ;
        RECT  1.480 -0.210 1.740 0.340 ;
        RECT  0.000 -0.210 1.480 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.225 2.310 8.400 2.730 ;
        RECT  8.055 1.845 8.225 2.730 ;
        RECT  7.505 2.310 8.055 2.730 ;
        RECT  7.335 1.845 7.505 2.730 ;
        RECT  6.785 2.310 7.335 2.730 ;
        RECT  6.615 1.800 6.785 2.730 ;
        RECT  6.065 2.310 6.615 2.730 ;
        RECT  5.895 1.845 6.065 2.730 ;
        RECT  5.345 2.310 5.895 2.730 ;
        RECT  5.175 1.845 5.345 2.730 ;
        RECT  4.630 2.310 5.175 2.730 ;
        RECT  4.095 1.800 4.630 2.730 ;
        RECT  3.540 2.310 4.095 2.730 ;
        RECT  3.370 1.800 3.540 2.730 ;
        RECT  2.820 2.310 3.370 2.730 ;
        RECT  2.650 1.780 2.820 2.730 ;
        RECT  2.125 2.310 2.650 2.730 ;
        RECT  1.865 2.020 2.125 2.730 ;
        RECT  1.335 2.310 1.865 2.730 ;
        RECT  1.165 2.005 1.335 2.730 ;
        RECT  0.000 2.310 1.165 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.400 2.520 ;
        LAYER M1 ;
        RECT  4.670 1.210 7.090 1.330 ;
        RECT  3.515 0.910 7.030 1.050 ;
        RECT  4.535 1.210 4.670 1.630 ;
        RECT  3.915 1.495 4.535 1.630 ;
        RECT  3.715 1.495 3.915 2.160 ;
        RECT  3.210 1.495 3.715 1.630 ;
        RECT  3.345 0.435 3.515 1.050 ;
        RECT  2.795 0.905 3.345 1.025 ;
        RECT  3.180 1.495 3.210 2.000 ;
        RECT  3.010 1.495 3.180 2.035 ;
        RECT  2.980 1.495 3.010 2.000 ;
        RECT  2.505 1.495 2.980 1.630 ;
        RECT  2.625 0.435 2.795 1.025 ;
        RECT  2.075 0.575 2.625 0.695 ;
        RECT  2.245 1.495 2.505 1.875 ;
        RECT  1.260 1.755 2.245 1.875 ;
        RECT  2.120 0.840 2.145 0.960 ;
        RECT  1.965 0.840 2.120 1.635 ;
        RECT  1.905 0.465 2.075 0.695 ;
        RECT  1.315 0.840 1.965 0.960 ;
        RECT  1.500 1.515 1.965 1.635 ;
        RECT  0.975 0.465 1.905 0.585 ;
        RECT  1.265 0.735 1.315 0.960 ;
        RECT  1.145 0.735 1.265 1.320 ;
        RECT  1.140 1.445 1.260 1.875 ;
        RECT  0.735 1.200 1.145 1.320 ;
        RECT  0.615 1.445 1.140 1.565 ;
        RECT  0.760 1.760 1.020 2.140 ;
        RECT  0.805 0.405 0.975 0.865 ;
        RECT  0.255 0.405 0.805 0.575 ;
        RECT  0.255 2.005 0.760 2.140 ;
        RECT  0.445 0.695 0.615 1.825 ;
        RECT  0.085 0.405 0.255 2.140 ;
    END
END TBUFX20AD
MACRO TBUFX2AD
    CLASS CORE ;
    FOREIGN TBUFX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.700 1.145 2.730 1.375 ;
        RECT  2.530 0.350 2.700 1.980 ;
        END
        AntennaDiffArea 0.341 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 0.980 0.525 1.150 ;
        RECT  0.070 0.980 0.210 1.375 ;
        END
        AntennaGateArea 0.1098 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.555 1.145 1.890 1.375 ;
        END
        AntennaGateArea 0.065 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.255 -0.210 2.800 0.210 ;
        RECT  1.965 -0.210 2.255 0.660 ;
        RECT  0.680 -0.210 1.965 0.210 ;
        RECT  0.510 -0.210 0.680 0.535 ;
        RECT  0.000 -0.210 0.510 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.340 2.310 2.800 2.730 ;
        RECT  2.170 1.550 2.340 2.730 ;
        RECT  1.770 1.685 2.170 1.805 ;
        RECT  0.275 2.310 2.170 2.730 ;
        RECT  0.105 1.740 0.275 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  1.840 0.855 2.135 1.025 ;
        RECT  1.435 2.020 2.050 2.140 ;
        RECT  1.720 0.390 1.840 1.025 ;
        RECT  1.700 0.390 1.720 0.510 ;
        RECT  1.440 0.350 1.700 0.510 ;
        RECT  1.435 0.690 1.535 0.950 ;
        RECT  1.175 0.390 1.440 0.510 ;
        RECT  1.315 0.690 1.435 2.140 ;
        RECT  0.690 2.020 1.315 2.140 ;
        RECT  1.055 0.390 1.175 1.775 ;
        RECT  0.835 0.390 1.055 0.535 ;
        RECT  0.850 1.655 1.055 1.775 ;
        RECT  0.810 0.675 0.930 1.410 ;
        RECT  0.295 0.675 0.810 0.800 ;
        RECT  0.640 1.270 0.810 1.410 ;
        RECT  0.450 1.880 0.690 2.140 ;
        RECT  0.520 1.270 0.640 1.735 ;
        RECT  0.125 0.365 0.295 0.800 ;
    END
END TBUFX2AD
MACRO TBUFX3AD
    CLASS CORE ;
    FOREIGN TBUFX3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.145 2.730 1.375 ;
        RECT  2.585 0.415 2.610 2.035 ;
        RECT  2.465 0.415 2.585 2.080 ;
        RECT  2.440 0.415 2.465 2.035 ;
        END
        AntennaDiffArea 0.318 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.045 0.560 1.375 ;
        RECT  0.130 1.045 0.350 1.215 ;
        END
        AntennaGateArea 0.1208 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.910 1.145 2.200 1.375 ;
        END
        AntennaGateArea 0.093 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 -0.210 3.080 0.210 ;
        RECT  2.800 -0.210 2.970 0.845 ;
        RECT  2.265 -0.210 2.800 0.210 ;
        RECT  2.045 -0.210 2.265 0.850 ;
        RECT  0.675 -0.210 2.045 0.210 ;
        RECT  0.505 -0.210 0.675 0.575 ;
        RECT  0.000 -0.210 0.505 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.970 2.310 3.080 2.730 ;
        RECT  2.800 1.590 2.970 2.730 ;
        RECT  2.240 2.310 2.800 2.730 ;
        RECT  2.070 1.510 2.240 2.730 ;
        RECT  0.265 2.310 2.070 2.730 ;
        RECT  0.095 1.520 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  1.695 0.390 1.865 0.905 ;
        RECT  1.505 1.525 1.865 1.695 ;
        RECT  1.470 1.960 1.700 2.190 ;
        RECT  1.195 0.390 1.695 0.510 ;
        RECT  1.470 0.735 1.505 1.695 ;
        RECT  1.440 0.735 1.470 2.190 ;
        RECT  1.325 0.735 1.440 2.130 ;
        RECT  0.485 1.960 1.325 2.130 ;
        RECT  1.075 0.390 1.195 1.740 ;
        RECT  0.890 0.390 1.075 0.575 ;
        RECT  0.815 0.710 0.935 1.675 ;
        RECT  0.280 0.710 0.815 0.830 ;
        RECT  0.440 1.500 0.815 1.675 ;
        RECT  0.110 0.405 0.280 0.830 ;
    END
END TBUFX3AD
MACRO TBUFX4AD
    CLASS CORE ;
    FOREIGN TBUFX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.385 0.375 2.575 2.085 ;
        RECT  2.310 0.725 2.385 1.235 ;
        END
        AntennaDiffArea 0.444 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 0.980 0.615 1.150 ;
        RECT  0.350 0.865 0.490 1.150 ;
        RECT  0.185 0.980 0.350 1.150 ;
        END
        AntennaGateArea 0.117 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.995 1.025 2.170 1.375 ;
        RECT  1.860 1.025 1.995 1.285 ;
        END
        AntennaGateArea 0.1137 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.985 -0.210 3.080 0.210 ;
        RECT  2.815 -0.210 2.985 0.890 ;
        RECT  2.190 -0.210 2.815 0.210 ;
        RECT  2.070 -0.210 2.190 0.840 ;
        RECT  0.635 -0.210 2.070 0.210 ;
        RECT  0.375 -0.210 0.635 0.255 ;
        RECT  0.000 -0.210 0.375 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.940 2.310 3.080 2.730 ;
        RECT  2.770 1.550 2.940 2.730 ;
        RECT  2.140 2.310 2.770 2.730 ;
        RECT  1.970 1.515 2.140 2.730 ;
        RECT  0.390 2.310 1.970 2.730 ;
        RECT  0.220 1.375 0.390 2.730 ;
        RECT  0.000 2.310 0.220 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  1.660 0.380 1.855 0.790 ;
        RECT  1.740 1.385 1.770 1.815 ;
        RECT  1.600 1.080 1.740 2.140 ;
        RECT  1.305 0.380 1.660 0.500 ;
        RECT  1.470 1.080 1.600 1.200 ;
        RECT  1.070 2.010 1.600 2.140 ;
        RECT  1.350 0.620 1.470 1.200 ;
        RECT  1.230 1.475 1.435 1.595 ;
        RECT  1.230 0.330 1.305 0.500 ;
        RECT  1.110 0.330 1.230 1.595 ;
        RECT  1.045 0.330 1.110 0.500 ;
        RECT  0.900 1.710 1.070 2.140 ;
        RECT  0.755 0.380 1.045 0.500 ;
        RECT  0.895 1.175 0.985 1.475 ;
        RECT  0.725 2.010 0.900 2.140 ;
        RECT  0.775 0.660 0.895 1.475 ;
        RECT  0.715 0.660 0.775 0.795 ;
        RECT  0.750 1.305 0.775 1.475 ;
        RECT  0.580 1.305 0.750 1.545 ;
        RECT  0.605 1.850 0.725 2.140 ;
        RECT  0.600 0.625 0.715 0.795 ;
        RECT  0.235 0.625 0.600 0.745 ;
        RECT  0.115 0.565 0.235 0.825 ;
    END
END TBUFX4AD
MACRO TBUFX6AD
    CLASS CORE ;
    FOREIGN TBUFX6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.645 0.385 3.815 2.065 ;
        RECT  3.095 1.095 3.645 1.375 ;
        RECT  2.925 0.445 3.095 2.070 ;
        RECT  2.870 0.585 2.925 1.375 ;
        END
        AntennaDiffArea 0.72 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.085 0.590 1.255 ;
        RECT  0.070 1.085 0.210 1.395 ;
        END
        AntennaGateArea 0.1173 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.145 2.170 1.400 ;
        RECT  1.715 1.230 2.030 1.400 ;
        END
        AntennaGateArea 0.192 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.455 -0.210 3.920 0.210 ;
        RECT  3.285 -0.210 3.455 0.770 ;
        RECT  2.725 -0.210 3.285 0.210 ;
        RECT  2.575 -0.210 2.725 0.810 ;
        RECT  2.145 -0.210 2.575 0.210 ;
        RECT  1.885 -0.210 2.145 0.250 ;
        RECT  0.690 -0.210 1.885 0.210 ;
        RECT  0.430 -0.210 0.690 0.510 ;
        RECT  0.000 -0.210 0.430 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.465 2.310 3.920 2.730 ;
        RECT  3.295 1.545 3.465 2.730 ;
        RECT  2.735 2.310 3.295 2.730 ;
        RECT  2.585 1.570 2.735 2.730 ;
        RECT  2.020 2.310 2.585 2.730 ;
        RECT  1.760 1.835 2.020 2.730 ;
        RECT  0.275 2.310 1.760 2.730 ;
        RECT  0.105 1.695 0.275 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  2.435 0.970 2.620 1.090 ;
        RECT  2.335 1.215 2.455 1.690 ;
        RECT  2.290 0.660 2.435 1.090 ;
        RECT  2.310 1.530 2.335 1.690 ;
        RECT  2.190 1.530 2.310 2.075 ;
        RECT  1.695 0.660 2.290 0.780 ;
        RECT  1.590 1.530 2.190 1.690 ;
        RECT  1.575 0.380 1.695 0.780 ;
        RECT  1.445 0.915 1.590 2.125 ;
        RECT  1.070 0.380 1.575 0.500 ;
        RECT  1.360 0.915 1.445 1.050 ;
        RECT  0.670 1.970 1.445 2.125 ;
        RECT  1.190 0.655 1.360 1.050 ;
        RECT  1.170 1.590 1.255 1.785 ;
        RECT  1.070 1.185 1.170 1.785 ;
        RECT  1.050 0.380 1.070 1.785 ;
        RECT  0.950 0.380 1.050 1.305 ;
        RECT  0.835 0.380 0.950 0.550 ;
        RECT  0.830 1.425 0.930 1.850 ;
        RECT  0.810 0.690 0.830 1.850 ;
        RECT  0.710 0.690 0.810 1.565 ;
        RECT  0.660 0.690 0.710 0.890 ;
        RECT  0.530 1.395 0.710 1.565 ;
        RECT  0.550 1.865 0.670 2.125 ;
        RECT  0.240 0.770 0.660 0.890 ;
        RECT  0.120 0.335 0.240 0.890 ;
    END
END TBUFX6AD
MACRO TBUFX8AD
    CLASS CORE ;
    FOREIGN TBUFX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.830 0.365 4.020 2.145 ;
        RECT  3.295 1.005 3.830 1.515 ;
        RECT  3.115 0.370 3.295 2.145 ;
        END
        AntennaDiffArea 0.778 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.085 0.610 1.205 ;
        RECT  0.070 1.085 0.210 1.375 ;
        END
        AntennaGateArea 0.1642 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.940 1.145 2.200 1.375 ;
        END
        AntennaGateArea 0.258 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.380 -0.210 4.480 0.210 ;
        RECT  4.225 -0.210 4.380 0.855 ;
        RECT  3.655 -0.210 4.225 0.210 ;
        RECT  3.485 -0.210 3.655 0.830 ;
        RECT  2.935 -0.210 3.485 0.210 ;
        RECT  2.765 -0.210 2.935 0.830 ;
        RECT  2.195 -0.210 2.765 0.210 ;
        RECT  2.025 -0.210 2.195 0.750 ;
        RECT  0.745 -0.210 2.025 0.210 ;
        RECT  0.485 -0.210 0.745 0.500 ;
        RECT  0.000 -0.210 0.485 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.375 2.310 4.480 2.730 ;
        RECT  4.205 1.620 4.375 2.730 ;
        RECT  3.645 2.310 4.205 2.730 ;
        RECT  3.475 1.695 3.645 2.730 ;
        RECT  2.925 2.310 3.475 2.730 ;
        RECT  2.755 1.645 2.925 2.730 ;
        RECT  2.145 2.310 2.755 2.730 ;
        RECT  1.945 1.895 2.145 2.730 ;
        RECT  0.265 2.310 1.945 2.730 ;
        RECT  0.810 1.710 1.070 1.895 ;
        RECT  0.265 1.710 0.810 1.855 ;
        RECT  0.095 1.635 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
        LAYER M1 ;
        RECT  2.560 0.950 2.720 1.080 ;
        RECT  2.610 1.280 2.680 1.400 ;
        RECT  2.490 1.280 2.610 1.725 ;
        RECT  2.460 0.400 2.560 1.080 ;
        RECT  2.415 1.280 2.490 2.095 ;
        RECT  2.390 0.400 2.460 1.050 ;
        RECT  2.320 1.605 2.415 2.095 ;
        RECT  1.835 0.875 2.390 0.995 ;
        RECT  1.745 1.605 2.320 1.725 ;
        RECT  1.665 0.400 1.835 0.995 ;
        RECT  1.620 1.145 1.745 2.140 ;
        RECT  1.180 0.400 1.665 0.540 ;
        RECT  1.475 1.145 1.620 1.265 ;
        RECT  0.690 2.020 1.620 2.140 ;
        RECT  1.300 0.660 1.475 1.265 ;
        RECT  1.240 1.385 1.410 1.710 ;
        RECT  1.180 1.385 1.240 1.555 ;
        RECT  1.060 0.400 1.180 1.555 ;
        RECT  0.900 0.400 1.060 0.520 ;
        RECT  0.820 0.740 0.940 1.590 ;
        RECT  0.360 0.740 0.820 0.865 ;
        RECT  0.475 1.420 0.820 1.590 ;
        RECT  0.430 1.975 0.690 2.140 ;
        RECT  0.190 0.430 0.360 0.865 ;
    END
END TBUFX8AD
MACRO TBUFXLAD
    CLASS CORE ;
    FOREIGN TBUFXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.380 2.450 2.105 ;
        RECT  2.170 0.380 2.310 0.500 ;
        RECT  2.260 1.845 2.310 2.105 ;
        END
        AntennaDiffArea 0.14 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.115 0.515 1.375 ;
        END
        AntennaGateArea 0.0888 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.905 1.025 2.075 1.240 ;
        RECT  1.890 1.115 1.905 1.240 ;
        RECT  1.750 1.115 1.890 1.375 ;
        END
        AntennaGateArea 0.0404 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.050 -0.210 2.520 0.210 ;
        RECT  1.790 -0.210 2.050 0.500 ;
        RECT  0.675 -0.210 1.790 0.210 ;
        RECT  0.415 -0.210 0.675 0.665 ;
        RECT  0.000 -0.210 0.415 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.090 2.310 2.520 2.730 ;
        RECT  1.830 1.810 2.090 2.730 ;
        RECT  0.265 2.310 1.830 2.730 ;
        RECT  0.095 1.565 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.520 2.520 ;
        LAYER M1 ;
        RECT  2.060 0.620 2.180 0.880 ;
        RECT  2.050 1.365 2.170 1.680 ;
        RECT  1.670 0.620 2.060 0.740 ;
        RECT  1.630 1.555 2.050 1.680 ;
        RECT  1.595 0.865 1.755 0.985 ;
        RECT  1.550 0.380 1.670 0.740 ;
        RECT  1.595 1.555 1.630 2.130 ;
        RECT  1.510 0.865 1.595 2.130 ;
        RECT  1.325 0.380 1.550 0.500 ;
        RECT  1.475 0.865 1.510 1.680 ;
        RECT  0.450 2.010 1.510 2.130 ;
        RECT  1.205 0.380 1.325 1.890 ;
        RECT  0.965 0.380 1.205 0.500 ;
        RECT  1.040 1.770 1.205 1.890 ;
        RECT  0.880 1.520 1.035 1.640 ;
        RECT  0.845 0.380 0.965 0.735 ;
        RECT  0.760 0.855 0.880 1.640 ;
        RECT  0.265 0.855 0.760 0.975 ;
        RECT  0.460 1.520 0.760 1.640 ;
        RECT  0.095 0.475 0.265 0.975 ;
    END
END TBUFXLAD
MACRO TIEHIAD
    CLASS CORE ;
    FOREIGN TIEHIAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.425 0.770 1.930 ;
        RECT  0.515 1.425 0.630 1.650 ;
        END
        AntennaDiffArea 0.094 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.325 -0.210 0.840 0.210 ;
        RECT  0.155 -0.210 0.325 0.905 ;
        RECT  0.000 -0.210 0.155 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.335 2.310 0.840 2.730 ;
        RECT  0.155 1.480 0.335 2.730 ;
        RECT  0.000 2.310 0.155 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 0.840 2.520 ;
        LAYER M1 ;
        RECT  0.515 0.735 0.685 1.225 ;
        RECT  0.395 1.055 0.515 1.225 ;
    END
END TIEHIAD
MACRO TIELOAD
    CLASS CORE ;
    FOREIGN TIELOAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.685 0.585 0.770 0.815 ;
        RECT  0.515 0.585 0.685 0.920 ;
        END
        AntennaDiffArea 0.075 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.325 -0.210 0.840 0.210 ;
        RECT  0.155 -0.210 0.325 0.860 ;
        RECT  0.000 -0.210 0.155 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.325 2.310 0.840 2.730 ;
        RECT  0.155 1.375 0.325 2.730 ;
        RECT  0.000 2.310 0.155 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 0.840 2.520 ;
        LAYER M1 ;
        RECT  0.515 1.055 0.685 1.545 ;
        RECT  0.275 1.055 0.515 1.225 ;
    END
END TIELOAD
MACRO TLATNCAX12AD
    CLASS CORE ;
    FOREIGN TLATNCAX12AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.670 0.380 9.910 1.955 ;
        RECT  6.825 0.380 9.670 0.670 ;
        RECT  9.440 1.125 9.670 1.955 ;
        RECT  9.385 1.370 9.440 1.955 ;
        RECT  9.215 1.370 9.385 2.125 ;
        RECT  8.250 1.370 9.215 1.770 ;
        RECT  7.950 1.370 8.250 2.120 ;
        RECT  6.970 1.370 7.950 1.770 ;
        RECT  6.775 1.370 6.970 2.085 ;
        RECT  6.655 0.380 6.825 0.550 ;
        END
        AntennaDiffArea 1.176 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.120 1.425 2.170 1.655 ;
        RECT  2.000 1.230 2.120 1.655 ;
        END
        AntennaGateArea 0.603 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.535 1.120 0.710 1.240 ;
        RECT  0.300 1.120 0.535 1.330 ;
        RECT  0.190 1.120 0.300 1.240 ;
        END
        AntennaGateArea 0.459 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.250 -0.210 10.080 0.210 ;
        RECT  8.990 -0.210 9.250 0.260 ;
        RECT  8.280 -0.210 8.990 0.210 ;
        RECT  8.020 -0.210 8.280 0.260 ;
        RECT  7.300 -0.210 8.020 0.210 ;
        RECT  7.040 -0.210 7.300 0.260 ;
        RECT  6.440 -0.210 7.040 0.210 ;
        RECT  6.180 -0.210 6.440 0.260 ;
        RECT  5.860 -0.210 6.180 0.210 ;
        RECT  5.600 -0.210 5.860 0.260 ;
        RECT  4.585 -0.210 5.600 0.210 ;
        RECT  4.325 -0.210 4.585 0.315 ;
        RECT  3.280 -0.210 4.325 0.210 ;
        RECT  3.020 -0.210 3.280 0.390 ;
        RECT  2.030 -0.210 3.020 0.210 ;
        RECT  1.770 -0.210 2.030 0.630 ;
        RECT  1.400 -0.210 1.770 0.210 ;
        RECT  1.140 -0.210 1.400 0.330 ;
        RECT  0.615 -0.210 1.140 0.210 ;
        RECT  0.445 -0.210 0.615 0.725 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.995 2.310 10.080 2.730 ;
        RECT  9.825 2.075 9.995 2.730 ;
        RECT  8.820 2.310 9.825 2.730 ;
        RECT  8.560 2.130 8.820 2.730 ;
        RECT  7.600 2.310 8.560 2.730 ;
        RECT  7.340 1.930 7.600 2.730 ;
        RECT  6.360 2.310 7.340 2.730 ;
        RECT  5.840 2.130 6.360 2.730 ;
        RECT  4.550 2.310 5.840 2.730 ;
        RECT  4.290 2.130 4.550 2.730 ;
        RECT  3.310 2.310 4.290 2.730 ;
        RECT  3.050 2.130 3.310 2.730 ;
        RECT  2.040 2.310 3.050 2.730 ;
        RECT  1.780 2.130 2.040 2.730 ;
        RECT  1.400 2.310 1.780 2.730 ;
        RECT  1.140 2.290 1.400 2.730 ;
        RECT  0.660 2.310 1.140 2.730 ;
        RECT  0.400 1.710 0.660 2.730 ;
        RECT  0.000 2.310 0.400 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 10.080 2.520 ;
        LAYER M1 ;
        RECT  9.305 0.790 9.550 0.910 ;
        RECT  9.185 0.790 9.305 1.200 ;
        RECT  6.460 1.080 9.185 1.200 ;
        RECT  6.705 0.840 9.060 0.960 ;
        RECT  6.585 0.745 6.705 0.960 ;
        RECT  6.535 0.745 6.585 0.865 ;
        RECT  6.415 0.380 6.535 0.865 ;
        RECT  6.340 1.000 6.460 2.010 ;
        RECT  5.500 0.380 6.415 0.500 ;
        RECT  5.530 1.890 6.340 2.010 ;
        RECT  6.100 0.645 6.220 1.565 ;
        RECT  6.025 0.645 6.100 0.815 ;
        RECT  5.740 1.395 6.100 1.565 ;
        RECT  5.500 0.950 5.980 1.070 ;
        RECT  5.620 1.210 5.740 1.565 ;
        RECT  5.270 1.890 5.530 2.180 ;
        RECT  5.380 0.380 5.500 1.770 ;
        RECT  2.390 0.510 5.380 0.630 ;
        RECT  2.400 1.650 5.380 1.770 ;
        RECT  1.880 1.890 5.270 2.010 ;
        RECT  5.140 0.750 5.260 1.490 ;
        RECT  1.640 0.750 5.140 0.870 ;
        RECT  3.790 1.370 5.140 1.490 ;
        RECT  4.895 0.990 5.015 1.250 ;
        RECT  4.085 0.990 4.895 1.110 ;
        RECT  3.825 0.990 4.085 1.170 ;
        RECT  2.520 0.990 3.825 1.110 ;
        RECT  3.530 1.340 3.790 1.490 ;
        RECT  2.830 1.370 3.530 1.490 ;
        RECT  2.570 1.330 2.830 1.490 ;
        RECT  2.260 0.990 2.520 1.170 ;
        RECT  1.880 0.990 2.260 1.110 ;
        RECT  1.760 0.990 1.880 2.010 ;
        RECT  0.950 1.890 1.760 2.010 ;
        RECT  1.520 0.610 1.640 1.760 ;
        RECT  1.440 0.610 1.520 0.870 ;
        RECT  1.440 1.500 1.520 1.760 ;
        RECT  0.950 1.035 1.400 1.300 ;
        RECT  0.830 0.350 0.950 2.010 ;
        RECT  0.230 0.855 0.830 0.975 ;
        RECT  0.230 1.465 0.830 1.585 ;
        RECT  0.110 0.350 0.230 0.975 ;
        RECT  0.110 1.465 0.230 2.010 ;
    END
END TLATNCAX12AD
MACRO TLATNCAX16AD
    CLASS CORE ;
    FOREIGN TLATNCAX16AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.185 0.380 12.425 1.955 ;
        RECT  8.095 0.380 12.185 0.670 ;
        RECT  11.855 1.170 12.185 1.955 ;
        RECT  11.685 1.170 11.855 2.125 ;
        RECT  11.480 1.170 11.685 1.955 ;
        RECT  10.635 1.455 11.480 1.955 ;
        RECT  10.465 1.455 10.635 2.155 ;
        RECT  9.415 1.455 10.465 1.955 ;
        RECT  9.245 1.455 9.415 2.160 ;
        RECT  8.195 1.455 9.245 1.955 ;
        RECT  8.025 1.455 8.195 2.145 ;
        RECT  7.905 0.380 8.095 0.550 ;
        END
        AntennaDiffArea 1.548 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.425 2.730 1.655 ;
        RECT  2.400 1.230 2.520 1.655 ;
        END
        AntennaGateArea 0.726 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.815 1.120 0.880 1.240 ;
        RECT  0.560 1.120 0.815 1.330 ;
        RECT  0.360 1.120 0.560 1.240 ;
        END
        AntennaGateArea 0.61 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  11.360 -0.210 12.600 0.210 ;
        RECT  11.100 -0.210 11.360 0.260 ;
        RECT  10.500 -0.210 11.100 0.210 ;
        RECT  10.240 -0.210 10.500 0.260 ;
        RECT  9.565 -0.210 10.240 0.210 ;
        RECT  9.305 -0.210 9.565 0.260 ;
        RECT  8.550 -0.210 9.305 0.210 ;
        RECT  8.290 -0.210 8.550 0.260 ;
        RECT  7.690 -0.210 8.290 0.210 ;
        RECT  7.430 -0.210 7.690 0.260 ;
        RECT  7.145 -0.210 7.430 0.210 ;
        RECT  6.885 -0.210 7.145 0.260 ;
        RECT  6.265 -0.210 6.885 0.210 ;
        RECT  6.005 -0.210 6.265 0.260 ;
        RECT  4.995 -0.210 6.005 0.210 ;
        RECT  4.735 -0.210 4.995 0.390 ;
        RECT  3.690 -0.210 4.735 0.210 ;
        RECT  3.430 -0.210 3.690 0.390 ;
        RECT  2.440 -0.210 3.430 0.210 ;
        RECT  2.180 -0.210 2.440 0.630 ;
        RECT  1.810 -0.210 2.180 0.210 ;
        RECT  1.550 -0.210 1.810 0.330 ;
        RECT  0.985 -0.210 1.550 0.210 ;
        RECT  0.815 -0.210 0.985 0.725 ;
        RECT  0.255 -0.210 0.815 0.210 ;
        RECT  0.085 -0.210 0.255 0.725 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.465 2.310 12.600 2.730 ;
        RECT  12.295 2.075 12.465 2.730 ;
        RECT  11.290 2.310 12.295 2.730 ;
        RECT  11.030 2.130 11.290 2.730 ;
        RECT  10.070 2.310 11.030 2.730 ;
        RECT  9.810 2.130 10.070 2.730 ;
        RECT  8.850 2.310 9.810 2.730 ;
        RECT  8.590 2.130 8.850 2.730 ;
        RECT  7.610 2.310 8.590 2.730 ;
        RECT  7.090 2.130 7.610 2.730 ;
        RECT  6.265 2.310 7.090 2.730 ;
        RECT  6.005 2.130 6.265 2.730 ;
        RECT  4.960 2.310 6.005 2.730 ;
        RECT  4.700 2.130 4.960 2.730 ;
        RECT  3.720 2.310 4.700 2.730 ;
        RECT  3.460 2.130 3.720 2.730 ;
        RECT  2.440 2.310 3.460 2.730 ;
        RECT  2.180 2.130 2.440 2.730 ;
        RECT  1.750 2.310 2.180 2.730 ;
        RECT  1.490 2.130 1.750 2.730 ;
        RECT  0.985 2.310 1.490 2.730 ;
        RECT  0.815 1.765 0.985 2.730 ;
        RECT  0.255 2.310 0.815 2.730 ;
        RECT  0.085 1.685 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 12.600 2.520 ;
        LAYER M1 ;
        RECT  11.665 0.930 12.030 1.050 ;
        RECT  11.510 0.840 11.665 1.050 ;
        RECT  7.955 0.840 11.510 0.960 ;
        RECT  7.710 1.140 11.205 1.260 ;
        RECT  7.835 0.745 7.955 0.960 ;
        RECT  7.785 0.745 7.835 0.865 ;
        RECT  7.665 0.380 7.785 0.865 ;
        RECT  7.590 1.000 7.710 2.010 ;
        RECT  6.750 0.380 7.665 0.500 ;
        RECT  6.780 1.890 7.590 2.010 ;
        RECT  7.350 0.620 7.470 1.565 ;
        RECT  7.210 0.620 7.350 0.740 ;
        RECT  6.990 1.395 7.350 1.565 ;
        RECT  7.110 0.880 7.230 1.140 ;
        RECT  6.750 0.950 7.110 1.070 ;
        RECT  6.870 1.210 6.990 1.565 ;
        RECT  6.520 1.890 6.780 2.180 ;
        RECT  6.630 0.380 6.750 1.770 ;
        RECT  2.800 0.510 6.630 0.630 ;
        RECT  2.850 1.650 6.630 1.770 ;
        RECT  2.280 1.890 6.520 2.010 ;
        RECT  6.390 0.750 6.510 1.480 ;
        RECT  2.040 0.750 6.390 0.870 ;
        RECT  2.980 1.360 6.390 1.480 ;
        RECT  5.235 0.990 5.495 1.190 ;
        RECT  4.495 0.990 5.235 1.110 ;
        RECT  4.235 0.990 4.495 1.190 ;
        RECT  2.920 0.990 4.235 1.110 ;
        RECT  2.660 0.990 2.920 1.190 ;
        RECT  2.280 0.990 2.660 1.110 ;
        RECT  2.160 0.990 2.280 2.010 ;
        RECT  1.320 1.890 2.160 2.010 ;
        RECT  1.920 0.610 2.040 1.760 ;
        RECT  1.850 0.610 1.920 0.870 ;
        RECT  1.320 1.035 1.800 1.300 ;
        RECT  1.200 0.350 1.320 2.010 ;
        RECT  0.600 0.855 1.200 0.975 ;
        RECT  0.625 1.465 1.200 1.585 ;
        RECT  0.450 1.465 0.625 1.965 ;
        RECT  0.480 0.350 0.600 0.975 ;
    END
END TLATNCAX16AD
MACRO TLATNCAX20AD
    CLASS CORE ;
    FOREIGN TLATNCAX20AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  14.950 0.380 15.510 2.010 ;
        RECT  9.510 0.380 14.950 0.680 ;
        RECT  14.665 1.170 14.950 2.010 ;
        RECT  14.565 1.170 14.665 2.120 ;
        RECT  14.495 1.430 14.565 2.120 ;
        RECT  13.385 1.430 14.495 2.010 ;
        RECT  13.215 1.430 13.385 2.150 ;
        RECT  12.145 1.430 13.215 2.010 ;
        RECT  11.975 1.430 12.145 2.125 ;
        RECT  10.885 1.430 11.975 2.010 ;
        RECT  10.715 1.430 10.885 2.150 ;
        RECT  9.635 1.430 10.715 2.010 ;
        RECT  9.465 1.430 9.635 2.150 ;
        END
        AntennaDiffArea 2.064 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.030 2.805 1.375 ;
        END
        AntennaGateArea 0.968 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.305 1.060 1.420 1.330 ;
        END
        AntennaGateArea 0.755 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  14.535 -0.210 15.680 0.210 ;
        RECT  14.275 -0.210 14.535 0.260 ;
        RECT  13.565 -0.210 14.275 0.210 ;
        RECT  13.305 -0.210 13.565 0.260 ;
        RECT  12.625 -0.210 13.305 0.210 ;
        RECT  12.105 -0.210 12.625 0.260 ;
        RECT  11.420 -0.210 12.105 0.210 ;
        RECT  10.900 -0.210 11.420 0.260 ;
        RECT  10.215 -0.210 10.900 0.210 ;
        RECT  9.955 -0.210 10.215 0.260 ;
        RECT  9.035 -0.210 9.955 0.210 ;
        RECT  8.515 -0.210 9.035 0.260 ;
        RECT  7.780 -0.210 8.515 0.210 ;
        RECT  7.520 -0.210 7.780 0.330 ;
        RECT  6.520 -0.210 7.520 0.210 ;
        RECT  6.260 -0.210 6.520 0.430 ;
        RECT  5.260 -0.210 6.260 0.210 ;
        RECT  5.000 -0.210 5.260 0.425 ;
        RECT  3.980 -0.210 5.000 0.210 ;
        RECT  3.720 -0.210 3.980 0.380 ;
        RECT  2.680 -0.210 3.720 0.210 ;
        RECT  1.900 -0.210 2.680 0.265 ;
        RECT  1.350 -0.210 1.900 0.210 ;
        RECT  1.180 -0.210 1.350 0.650 ;
        RECT  0.630 -0.210 1.180 0.210 ;
        RECT  0.460 -0.210 0.630 0.650 ;
        RECT  0.000 -0.210 0.460 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.320 2.310 15.680 2.730 ;
        RECT  15.060 2.130 15.320 2.730 ;
        RECT  14.100 2.310 15.060 2.730 ;
        RECT  13.840 2.130 14.100 2.730 ;
        RECT  12.820 2.310 13.840 2.730 ;
        RECT  12.560 2.130 12.820 2.730 ;
        RECT  11.560 2.310 12.560 2.730 ;
        RECT  11.300 2.130 11.560 2.730 ;
        RECT  10.310 2.310 11.300 2.730 ;
        RECT  10.050 2.130 10.310 2.730 ;
        RECT  8.920 2.310 10.050 2.730 ;
        RECT  8.400 2.130 8.920 2.730 ;
        RECT  7.700 2.310 8.400 2.730 ;
        RECT  7.440 2.130 7.700 2.730 ;
        RECT  6.480 2.310 7.440 2.730 ;
        RECT  6.220 2.130 6.480 2.730 ;
        RECT  5.220 2.310 6.220 2.730 ;
        RECT  4.960 2.130 5.220 2.730 ;
        RECT  4.000 2.310 4.960 2.730 ;
        RECT  3.740 2.130 4.000 2.730 ;
        RECT  2.675 2.310 3.740 2.730 ;
        RECT  1.895 2.270 2.675 2.730 ;
        RECT  1.350 2.310 1.895 2.730 ;
        RECT  1.180 1.760 1.350 2.730 ;
        RECT  0.630 2.310 1.180 2.730 ;
        RECT  0.460 1.760 0.630 2.730 ;
        RECT  0.000 2.310 0.460 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 15.680 2.520 ;
        LAYER M1 ;
        RECT  14.445 0.900 14.830 1.020 ;
        RECT  14.325 0.900 14.445 1.260 ;
        RECT  9.150 1.140 14.325 1.260 ;
        RECT  9.390 0.850 14.205 0.970 ;
        RECT  9.270 0.380 9.390 0.970 ;
        RECT  8.070 0.380 9.270 0.500 ;
        RECT  9.030 1.040 9.150 2.010 ;
        RECT  8.110 1.890 9.030 2.010 ;
        RECT  8.790 0.645 8.910 1.480 ;
        RECT  8.735 0.645 8.790 0.815 ;
        RECT  8.715 1.360 8.790 1.480 ;
        RECT  8.545 1.360 8.715 1.575 ;
        RECT  8.550 0.960 8.670 1.220 ;
        RECT  8.070 1.010 8.550 1.130 ;
        RECT  8.190 1.360 8.545 1.480 ;
        RECT  7.850 1.890 8.110 2.190 ;
        RECT  7.950 0.380 8.070 1.770 ;
        RECT  7.840 0.550 7.950 0.860 ;
        RECT  3.345 1.650 7.950 1.770 ;
        RECT  2.815 1.890 7.850 2.010 ;
        RECT  3.090 0.550 7.840 0.670 ;
        RECT  7.590 1.070 7.830 1.330 ;
        RECT  7.470 0.790 7.590 1.480 ;
        RECT  2.470 0.790 7.470 0.910 ;
        RECT  3.240 1.360 7.470 1.480 ;
        RECT  3.045 1.070 7.270 1.190 ;
        RECT  3.175 1.600 3.345 1.770 ;
        RECT  2.925 1.070 3.045 1.620 ;
        RECT  2.815 1.495 2.925 1.620 ;
        RECT  2.695 1.495 2.815 2.010 ;
        RECT  1.710 1.805 2.695 1.925 ;
        RECT  2.350 0.665 2.470 1.685 ;
        RECT  2.210 0.665 2.350 0.910 ;
        RECT  2.210 1.515 2.350 1.685 ;
        RECT  1.710 1.070 2.230 1.190 ;
        RECT  1.540 0.435 1.710 1.925 ;
        RECT  0.990 0.770 1.540 0.890 ;
        RECT  0.990 1.520 1.540 1.640 ;
        RECT  0.820 0.435 0.990 0.890 ;
        RECT  0.820 1.520 0.990 1.950 ;
        RECT  0.270 0.770 0.820 0.890 ;
        RECT  0.270 1.520 0.820 1.640 ;
        RECT  0.100 0.430 0.270 0.890 ;
        RECT  0.100 1.520 0.270 1.950 ;
    END
END TLATNCAX20AD
MACRO TLATNCAX2AD
    CLASS CORE ;
    FOREIGN TLATNCAX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.545 1.425 3.570 1.655 ;
        RECT  3.375 1.425 3.545 2.035 ;
        RECT  3.265 1.425 3.375 1.655 ;
        RECT  3.140 0.680 3.265 1.655 ;
        RECT  3.015 0.680 3.140 0.850 ;
        END
        AntennaDiffArea 0.276 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.090 0.910 1.375 1.330 ;
        END
        AntennaGateArea 0.132 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.165 1.020 0.285 1.655 ;
        RECT  0.070 1.410 0.165 1.655 ;
        END
        AntennaGateArea 0.114 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.545 -0.210 3.640 0.210 ;
        RECT  3.425 -0.210 3.545 0.900 ;
        RECT  2.810 -0.210 3.425 0.210 ;
        RECT  3.385 0.640 3.425 0.900 ;
        RECT  2.290 -0.210 2.810 0.265 ;
        RECT  1.290 -0.210 2.290 0.210 ;
        RECT  1.030 -0.210 1.290 0.490 ;
        RECT  0.255 -0.210 1.030 0.210 ;
        RECT  0.085 -0.210 0.255 0.765 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.765 2.310 3.640 2.730 ;
        RECT  2.245 2.260 2.765 2.730 ;
        RECT  1.145 2.310 2.245 2.730 ;
        RECT  0.885 2.130 1.145 2.730 ;
        RECT  0.315 2.310 0.885 2.730 ;
        RECT  0.145 2.265 0.315 2.730 ;
        RECT  0.000 2.310 0.145 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  3.135 0.330 3.305 0.550 ;
        RECT  2.780 0.430 3.135 0.550 ;
        RECT  2.900 1.035 3.020 2.140 ;
        RECT  1.385 2.020 2.900 2.140 ;
        RECT  2.660 0.430 2.780 1.900 ;
        RECT  2.160 0.430 2.660 0.550 ;
        RECT  2.580 1.120 2.660 1.380 ;
        RECT  1.520 1.780 2.660 1.900 ;
        RECT  2.460 1.500 2.540 1.660 ;
        RECT  2.460 0.705 2.485 0.875 ;
        RECT  2.280 0.705 2.460 1.660 ;
        RECT  2.170 1.120 2.280 1.380 ;
        RECT  2.040 0.370 2.160 0.550 ;
        RECT  1.640 0.370 2.040 0.490 ;
        RECT  1.920 0.795 1.980 1.315 ;
        RECT  1.680 1.520 1.970 1.640 ;
        RECT  1.800 0.610 1.920 1.315 ;
        RECT  0.940 0.610 1.800 0.730 ;
        RECT  1.535 0.850 1.680 1.640 ;
        RECT  1.385 1.520 1.535 1.640 ;
        RECT  1.265 1.520 1.385 2.140 ;
        RECT  0.525 1.890 1.265 2.010 ;
        RECT  0.885 0.610 0.940 1.710 ;
        RECT  0.820 0.345 0.885 1.710 ;
        RECT  0.750 0.345 0.820 0.730 ;
        RECT  0.665 1.450 0.820 1.710 ;
        RECT  0.715 0.345 0.750 0.515 ;
        RECT  0.590 0.985 0.700 1.245 ;
        RECT  0.525 0.670 0.590 1.245 ;
        RECT  0.520 0.670 0.525 2.010 ;
        RECT  0.405 0.670 0.520 2.050 ;
        RECT  0.345 1.790 0.405 2.050 ;
    END
END TLATNCAX2AD
MACRO TLATNCAX3AD
    CLASS CORE ;
    FOREIGN TLATNCAX3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.200 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.410 0.660 3.660 0.780 ;
        RECT  3.505 1.285 3.570 1.795 ;
        RECT  3.410 1.285 3.505 1.865 ;
        RECT  3.335 0.660 3.410 1.865 ;
        RECT  3.290 0.660 3.335 1.435 ;
        END
        AntennaDiffArea 0.282 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.020 1.330 1.655 ;
        END
        AntennaGateArea 0.15 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.160 1.005 0.305 1.375 ;
        RECT  0.070 1.145 0.160 1.375 ;
        END
        AntennaGateArea 0.137 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.050 -0.210 4.200 0.210 ;
        RECT  3.790 -0.210 4.050 0.300 ;
        RECT  3.280 -0.210 3.790 0.210 ;
        RECT  3.020 -0.210 3.280 0.300 ;
        RECT  2.560 -0.210 3.020 0.210 ;
        RECT  2.300 -0.210 2.560 0.300 ;
        RECT  1.240 -0.210 2.300 0.210 ;
        RECT  0.980 -0.210 1.240 0.390 ;
        RECT  0.680 -0.210 0.980 0.210 ;
        RECT  0.420 -0.210 0.680 0.450 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.090 2.310 4.200 2.730 ;
        RECT  3.970 1.540 4.090 2.730 ;
        RECT  2.910 2.310 3.970 2.730 ;
        RECT  2.390 2.210 2.910 2.730 ;
        RECT  1.160 2.310 2.390 2.730 ;
        RECT  0.900 2.210 1.160 2.730 ;
        RECT  0.680 2.310 0.900 2.730 ;
        RECT  0.420 2.210 0.680 2.730 ;
        RECT  0.000 2.310 0.420 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.200 2.520 ;
        LAYER M1 ;
        RECT  3.850 1.200 4.115 1.320 ;
        RECT  3.780 0.420 3.900 1.060 ;
        RECT  3.730 1.200 3.850 2.105 ;
        RECT  2.300 0.420 3.780 0.540 ;
        RECT  3.530 0.940 3.780 1.060 ;
        RECT  3.120 1.985 3.730 2.105 ;
        RECT  3.000 0.890 3.120 2.105 ;
        RECT  2.080 1.930 3.000 2.050 ;
        RECT  2.760 0.660 2.880 1.750 ;
        RECT  2.620 0.660 2.760 0.780 ;
        RECT  2.375 1.630 2.760 1.750 ;
        RECT  2.520 1.000 2.640 1.260 ;
        RECT  2.300 1.000 2.520 1.175 ;
        RECT  2.255 1.340 2.375 1.750 ;
        RECT  2.180 0.420 2.300 1.175 ;
        RECT  2.115 1.340 2.255 1.500 ;
        RECT  1.630 0.420 2.180 0.540 ;
        RECT  1.995 1.055 2.180 1.175 ;
        RECT  1.960 1.620 2.080 2.050 ;
        RECT  1.870 0.660 2.020 0.920 ;
        RECT  1.875 1.055 1.995 1.400 ;
        RECT  1.570 1.930 1.960 2.050 ;
        RECT  1.820 1.280 1.875 1.400 ;
        RECT  0.925 0.660 1.870 0.780 ;
        RECT  1.700 1.280 1.820 1.810 ;
        RECT  1.570 0.980 1.730 1.100 ;
        RECT  1.450 0.980 1.570 2.050 ;
        RECT  0.230 1.930 1.450 2.050 ;
        RECT  0.805 0.660 0.925 1.595 ;
        RECT  0.755 0.660 0.805 0.905 ;
        RECT  0.755 1.425 0.805 1.595 ;
        RECT  0.610 1.000 0.680 1.260 ;
        RECT  0.490 0.765 0.610 1.620 ;
        RECT  0.230 0.765 0.490 0.885 ;
        RECT  0.230 1.500 0.490 1.620 ;
        RECT  0.110 0.550 0.230 0.885 ;
        RECT  0.110 1.500 0.230 2.050 ;
    END
END TLATNCAX3AD
MACRO TLATNCAX4AD
    CLASS CORE ;
    FOREIGN TLATNCAX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.360 0.490 5.490 1.610 ;
        RECT  4.610 0.490 5.360 0.620 ;
        RECT  4.805 1.450 5.360 1.610 ;
        RECT  4.625 1.450 4.805 2.015 ;
        END
        AntennaDiffArea 0.38 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.690 0.990 2.730 1.375 ;
        RECT  2.570 0.990 2.690 1.590 ;
        RECT  1.455 1.470 2.570 1.590 ;
        RECT  1.285 1.135 1.455 1.590 ;
        END
        AntennaGateArea 0.226 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.230 1.085 0.375 1.255 ;
        RECT  0.070 1.085 0.230 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.260 -0.210 5.600 0.210 ;
        RECT  5.000 -0.210 5.260 0.310 ;
        RECT  4.460 -0.210 5.000 0.210 ;
        RECT  4.300 -0.210 4.460 0.700 ;
        RECT  2.930 -0.210 4.300 0.210 ;
        RECT  2.670 -0.210 2.930 0.260 ;
        RECT  1.360 -0.210 2.670 0.210 ;
        RECT  1.100 -0.210 1.360 0.280 ;
        RECT  0.255 -0.210 1.100 0.210 ;
        RECT  0.085 -0.210 0.255 0.830 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.415 2.310 5.600 2.730 ;
        RECT  5.245 1.755 5.415 2.730 ;
        RECT  4.170 2.310 5.245 2.730 ;
        RECT  3.390 2.210 4.170 2.730 ;
        RECT  2.625 2.310 3.390 2.730 ;
        RECT  2.365 2.210 2.625 2.730 ;
        RECT  1.340 2.310 2.365 2.730 ;
        RECT  1.080 2.210 1.340 2.730 ;
        RECT  0.255 2.310 1.080 2.730 ;
        RECT  0.085 1.540 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  5.120 0.960 5.240 1.220 ;
        RECT  4.180 1.100 5.120 1.220 ;
        RECT  4.180 0.860 4.730 0.980 ;
        RECT  4.060 0.380 4.180 0.980 ;
        RECT  4.060 1.100 4.180 2.015 ;
        RECT  3.700 0.380 4.060 0.500 ;
        RECT  3.275 1.895 4.060 2.015 ;
        RECT  3.820 0.620 3.940 1.600 ;
        RECT  3.360 1.480 3.820 1.600 ;
        RECT  3.580 0.380 3.700 1.280 ;
        RECT  1.730 0.415 3.580 0.535 ;
        RECT  2.970 1.080 3.580 1.200 ;
        RECT  3.240 1.340 3.360 1.600 ;
        RECT  3.200 0.675 3.340 0.935 ;
        RECT  3.155 1.895 3.275 2.090 ;
        RECT  2.450 0.675 3.200 0.795 ;
        RECT  3.090 1.970 3.155 2.090 ;
        RECT  2.830 1.970 3.090 2.190 ;
        RECT  2.850 1.080 2.970 1.850 ;
        RECT  1.730 1.730 2.850 1.850 ;
        RECT  0.635 1.970 2.830 2.090 ;
        RECT  2.330 0.675 2.450 1.350 ;
        RECT  1.870 1.230 2.330 1.350 ;
        RECT  2.030 0.950 2.210 1.070 ;
        RECT  1.910 0.655 2.030 1.070 ;
        RECT  1.505 0.655 1.910 0.775 ;
        RECT  1.730 1.190 1.870 1.350 ;
        RECT  1.610 0.895 1.730 1.350 ;
        RECT  1.130 0.895 1.610 1.015 ;
        RECT  1.385 0.410 1.505 0.775 ;
        RECT  0.635 0.410 1.385 0.530 ;
        RECT  1.010 0.670 1.130 1.695 ;
        RECT  0.760 0.670 1.010 0.790 ;
        RECT  0.805 1.525 1.010 1.695 ;
        RECT  0.635 0.985 0.890 1.245 ;
        RECT  0.515 0.410 0.635 2.090 ;
        RECT  0.445 0.410 0.515 0.840 ;
        RECT  0.470 1.455 0.515 2.090 ;
    END
END TLATNCAX4AD
MACRO TLATNCAX6AD
    CLASS CORE ;
    FOREIGN TLATNCAX6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.160 0.435 6.340 2.030 ;
        RECT  6.150 0.435 6.160 1.610 ;
        RECT  4.890 0.435 6.150 0.625 ;
        RECT  5.090 1.420 6.150 1.610 ;
        RECT  4.900 1.420 5.090 2.060 ;
        END
        AntennaDiffArea 0.664 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 0.990 3.010 1.375 ;
        RECT  2.850 0.990 2.970 1.610 ;
        RECT  1.740 1.490 2.850 1.610 ;
        RECT  1.620 1.135 1.740 1.610 ;
        RECT  1.565 1.135 1.620 1.305 ;
        END
        AntennaGateArea 0.3 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.290 1.110 0.550 1.375 ;
        END
        AntennaGateArea 0.24 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.320 -0.210 6.440 0.210 ;
        RECT  6.060 -0.210 6.320 0.310 ;
        RECT  5.540 -0.210 6.060 0.210 ;
        RECT  5.280 -0.210 5.540 0.310 ;
        RECT  4.740 -0.210 5.280 0.210 ;
        RECT  4.580 -0.210 4.740 0.700 ;
        RECT  3.210 -0.210 4.580 0.210 ;
        RECT  2.950 -0.210 3.210 0.260 ;
        RECT  1.590 -0.210 2.950 0.210 ;
        RECT  0.810 -0.210 1.590 0.280 ;
        RECT  0.255 -0.210 0.810 0.210 ;
        RECT  0.085 -0.210 0.255 0.885 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 2.310 6.440 2.730 ;
        RECT  5.545 1.730 5.715 2.730 ;
        RECT  4.450 2.310 5.545 2.730 ;
        RECT  3.670 2.210 4.450 2.730 ;
        RECT  2.950 2.310 3.670 2.730 ;
        RECT  2.690 2.210 2.950 2.730 ;
        RECT  1.590 2.310 2.690 2.730 ;
        RECT  0.810 2.210 1.590 2.730 ;
        RECT  0.260 2.310 0.810 2.730 ;
        RECT  0.100 1.500 0.260 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.440 2.520 ;
        LAYER M1 ;
        RECT  5.910 0.800 6.030 1.060 ;
        RECT  5.010 0.840 5.910 0.960 ;
        RECT  4.460 1.100 5.620 1.220 ;
        RECT  4.750 0.840 5.010 0.980 ;
        RECT  4.460 0.840 4.750 0.960 ;
        RECT  4.340 0.380 4.460 0.960 ;
        RECT  4.340 1.100 4.460 2.015 ;
        RECT  3.980 0.380 4.340 0.500 ;
        RECT  3.555 1.895 4.340 2.015 ;
        RECT  4.100 0.620 4.220 1.600 ;
        RECT  3.640 1.480 4.100 1.600 ;
        RECT  3.860 0.380 3.980 1.280 ;
        RECT  2.010 0.415 3.860 0.535 ;
        RECT  3.250 1.080 3.860 1.200 ;
        RECT  3.520 1.340 3.640 1.600 ;
        RECT  3.480 0.675 3.620 0.935 ;
        RECT  3.435 1.895 3.555 2.090 ;
        RECT  2.730 0.675 3.480 0.795 ;
        RECT  3.370 1.970 3.435 2.090 ;
        RECT  3.110 1.970 3.370 2.190 ;
        RECT  3.130 1.080 3.250 1.850 ;
        RECT  2.010 1.730 3.130 1.850 ;
        RECT  1.755 1.970 3.110 2.090 ;
        RECT  2.610 0.675 2.730 1.350 ;
        RECT  2.150 1.230 2.610 1.350 ;
        RECT  2.310 0.950 2.490 1.070 ;
        RECT  2.190 0.655 2.310 1.070 ;
        RECT  1.785 0.655 2.190 0.775 ;
        RECT  2.010 1.190 2.150 1.350 ;
        RECT  1.890 0.895 2.010 1.350 ;
        RECT  1.410 0.895 1.890 1.015 ;
        RECT  1.665 0.450 1.785 0.775 ;
        RECT  1.635 1.895 1.755 2.090 ;
        RECT  0.590 0.450 1.665 0.570 ;
        RECT  0.790 1.895 1.635 2.015 ;
        RECT  1.290 0.690 1.410 1.710 ;
        RECT  1.040 0.690 1.290 0.810 ;
        RECT  1.085 1.540 1.290 1.710 ;
        RECT  1.050 0.985 1.170 1.245 ;
        RECT  0.790 0.985 1.050 1.105 ;
        RECT  0.670 0.870 0.790 2.015 ;
        RECT  0.590 0.870 0.670 0.990 ;
        RECT  0.470 1.495 0.670 2.015 ;
        RECT  0.470 0.450 0.590 0.990 ;
    END
END TLATNCAX6AD
MACRO TLATNCAX8AD
    CLASS CORE ;
    FOREIGN TLATNCAX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.560 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.270 0.435 7.460 1.610 ;
        RECT  5.450 0.435 7.270 0.625 ;
        RECT  7.120 1.420 7.270 1.610 ;
        RECT  6.540 1.420 7.120 2.030 ;
        RECT  5.650 1.420 6.540 1.705 ;
        RECT  5.460 1.420 5.650 2.060 ;
        END
        AntennaDiffArea 0.764 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.425 0.990 3.570 1.610 ;
        RECT  2.330 1.490 3.425 1.610 ;
        RECT  2.180 1.190 2.330 1.610 ;
        RECT  2.070 1.190 2.180 1.310 ;
        END
        AntennaGateArea 0.414 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.290 1.120 0.550 1.375 ;
        END
        AntennaGateArea 0.312 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.880 -0.210 7.560 0.210 ;
        RECT  6.620 -0.210 6.880 0.310 ;
        RECT  6.100 -0.210 6.620 0.210 ;
        RECT  5.840 -0.210 6.100 0.310 ;
        RECT  5.300 -0.210 5.840 0.210 ;
        RECT  5.140 -0.210 5.300 0.700 ;
        RECT  3.770 -0.210 5.140 0.210 ;
        RECT  3.510 -0.210 3.770 0.260 ;
        RECT  2.465 -0.210 3.510 0.210 ;
        RECT  2.205 -0.210 2.465 0.295 ;
        RECT  1.040 -0.210 2.205 0.210 ;
        RECT  0.780 -0.210 1.040 0.280 ;
        RECT  0.255 -0.210 0.780 0.210 ;
        RECT  0.085 -0.210 0.255 0.885 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.475 2.310 7.560 2.730 ;
        RECT  7.305 1.730 7.475 2.730 ;
        RECT  6.255 2.310 7.305 2.730 ;
        RECT  6.085 2.035 6.255 2.730 ;
        RECT  5.010 2.310 6.085 2.730 ;
        RECT  4.230 2.210 5.010 2.730 ;
        RECT  3.490 2.310 4.230 2.730 ;
        RECT  3.230 2.210 3.490 2.730 ;
        RECT  2.230 2.310 3.230 2.730 ;
        RECT  1.970 2.210 2.230 2.730 ;
        RECT  1.015 2.310 1.970 2.730 ;
        RECT  0.845 2.150 1.015 2.730 ;
        RECT  0.255 2.310 0.845 2.730 ;
        RECT  0.085 1.560 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.560 2.520 ;
        LAYER M1 ;
        RECT  6.815 0.780 6.935 1.220 ;
        RECT  5.020 1.100 6.815 1.220 ;
        RECT  5.020 0.860 6.670 0.980 ;
        RECT  4.900 0.380 5.020 0.980 ;
        RECT  4.900 1.100 5.020 2.015 ;
        RECT  4.540 0.380 4.900 0.500 ;
        RECT  4.050 1.895 4.900 2.015 ;
        RECT  4.660 0.620 4.780 1.600 ;
        RECT  4.200 1.480 4.660 1.600 ;
        RECT  4.420 0.380 4.540 1.280 ;
        RECT  1.765 0.415 4.420 0.535 ;
        RECT  3.810 1.080 4.420 1.200 ;
        RECT  4.080 1.340 4.200 1.600 ;
        RECT  4.040 0.675 4.180 0.935 ;
        RECT  3.930 1.895 4.050 2.130 ;
        RECT  3.305 0.675 4.040 0.795 ;
        RECT  3.670 1.970 3.930 2.130 ;
        RECT  3.690 1.080 3.810 1.850 ;
        RECT  1.555 1.730 3.690 1.850 ;
        RECT  1.815 1.970 3.670 2.090 ;
        RECT  3.185 0.675 3.305 1.350 ;
        RECT  2.730 1.230 3.185 1.350 ;
        RECT  2.870 0.950 3.065 1.070 ;
        RECT  2.750 0.710 2.870 1.070 ;
        RECT  1.525 0.710 2.750 0.830 ;
        RECT  2.570 1.190 2.730 1.350 ;
        RECT  2.450 0.950 2.570 1.350 ;
        RECT  1.720 0.950 2.450 1.070 ;
        RECT  1.690 1.970 1.815 2.140 ;
        RECT  1.645 0.330 1.765 0.590 ;
        RECT  1.460 0.950 1.720 1.310 ;
        RECT  1.260 2.020 1.690 2.140 ;
        RECT  1.385 1.730 1.555 1.900 ;
        RECT  1.405 0.450 1.525 0.830 ;
        RECT  1.285 0.950 1.460 1.070 ;
        RECT  0.590 0.450 1.405 0.570 ;
        RECT  1.160 0.725 1.285 1.545 ;
        RECT  1.140 1.835 1.260 2.140 ;
        RECT  1.115 0.725 1.160 0.905 ;
        RECT  1.115 1.375 1.160 1.545 ;
        RECT  0.955 1.835 1.140 1.955 ;
        RECT  0.955 1.015 1.040 1.275 ;
        RECT  0.835 0.870 0.955 1.955 ;
        RECT  0.590 0.870 0.835 0.990 ;
        RECT  0.615 1.835 0.835 1.955 ;
        RECT  0.445 1.525 0.615 1.955 ;
        RECT  0.470 0.450 0.590 0.990 ;
    END
END TLATNCAX8AD
MACRO TLATNSRX1AD
    CLASS CORE ;
    FOREIGN TLATNSRX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.880 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.065 0.230 1.325 ;
        RECT  0.070 1.065 0.210 1.655 ;
        END
        AntennaGateArea 0.074 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.865 1.960 1.330 ;
        END
        AntennaGateArea 0.124 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.670 0.495 5.810 1.920 ;
        RECT  5.640 0.495 5.670 0.755 ;
        RECT  5.640 1.400 5.670 1.920 ;
        END
        AntennaDiffArea 0.209 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.985 0.540 5.075 0.710 ;
        RECT  4.985 1.390 5.035 1.820 ;
        RECT  4.865 0.540 4.985 1.820 ;
        RECT  4.830 0.865 4.865 1.375 ;
        END
        AntennaDiffArea 0.209 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.980 0.745 4.170 1.095 ;
        END
        AntennaGateArea 0.068 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.420 0.865 1.610 1.325 ;
        END
        AntennaGateArea 0.123 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.430 -0.210 5.880 0.210 ;
        RECT  5.270 -0.210 5.430 0.745 ;
        RECT  4.360 -0.210 5.270 0.210 ;
        RECT  4.180 -0.210 4.360 0.620 ;
        RECT  3.300 -0.210 4.180 0.210 ;
        RECT  3.040 -0.210 3.300 0.345 ;
        RECT  1.425 -0.210 3.040 0.210 ;
        RECT  1.255 -0.210 1.425 0.430 ;
        RECT  0.230 -0.210 1.255 0.210 ;
        RECT  0.070 -0.210 0.230 0.830 ;
        RECT  0.000 -0.210 0.070 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.460 2.310 5.880 2.730 ;
        RECT  5.200 2.220 5.460 2.730 ;
        RECT  4.360 2.310 5.200 2.730 ;
        RECT  4.100 2.220 4.360 2.730 ;
        RECT  3.340 2.310 4.100 2.730 ;
        RECT  3.080 2.015 3.340 2.730 ;
        RECT  1.810 2.310 3.080 2.730 ;
        RECT  1.550 2.220 1.810 2.730 ;
        RECT  0.230 2.310 1.550 2.730 ;
        RECT  0.070 1.775 0.230 2.730 ;
        RECT  0.000 2.310 0.070 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.880 2.520 ;
        LAYER M1 ;
        RECT  5.480 1.015 5.530 1.275 ;
        RECT  5.360 1.015 5.480 2.100 ;
        RECT  4.710 1.980 5.360 2.100 ;
        RECT  4.590 0.450 4.710 2.100 ;
        RECT  4.530 0.450 4.590 0.710 ;
        RECT  4.550 1.650 4.590 2.100 ;
        RECT  3.850 1.980 4.550 2.100 ;
        RECT  4.410 1.010 4.470 1.270 ;
        RECT  4.290 1.010 4.410 1.860 ;
        RECT  0.930 1.740 4.290 1.860 ;
        RECT  3.860 0.455 3.975 0.625 ;
        RECT  3.860 1.215 3.950 1.600 ;
        RECT  3.830 0.455 3.860 1.600 ;
        RECT  3.590 1.980 3.850 2.190 ;
        RECT  3.740 0.455 3.830 1.335 ;
        RECT  3.470 1.215 3.740 1.335 ;
        RECT  2.200 1.500 3.680 1.620 ;
        RECT  3.490 0.495 3.610 1.005 ;
        RECT  2.200 0.885 3.490 1.005 ;
        RECT  3.210 1.150 3.470 1.335 ;
        RECT  2.320 1.215 3.210 1.335 ;
        RECT  2.400 1.980 2.660 2.190 ;
        RECT  0.590 1.980 2.400 2.100 ;
        RECT  1.020 0.550 2.390 0.670 ;
        RECT  2.080 0.885 2.200 1.620 ;
        RECT  1.170 1.500 2.080 1.620 ;
        RECT  1.050 1.120 1.170 1.620 ;
        RECT  0.860 1.120 1.050 1.380 ;
        RECT  0.900 0.550 1.020 1.000 ;
        RECT  0.810 1.500 0.930 1.860 ;
        RECT  0.710 0.880 0.900 1.000 ;
        RECT  0.680 0.330 0.820 0.450 ;
        RECT  0.710 1.500 0.810 1.620 ;
        RECT  0.590 0.880 0.710 1.620 ;
        RECT  0.560 0.330 0.680 0.760 ;
        RECT  0.470 1.780 0.590 2.100 ;
        RECT  0.470 0.640 0.560 0.760 ;
        RECT  0.350 0.640 0.470 1.900 ;
    END
END TLATNSRX1AD
MACRO TLATNSRX2AD
    CLASS CORE ;
    FOREIGN TLATNSRX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.230 1.375 ;
        END
        AntennaGateArea 0.091 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.070 1.990 1.375 ;
        RECT  1.750 0.865 1.890 1.375 ;
        END
        AntennaGateArea 0.152 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.950 0.365 6.090 2.045 ;
        RECT  5.920 0.365 5.950 0.885 ;
        RECT  5.920 1.525 5.950 2.045 ;
        END
        AntennaDiffArea 0.373 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 0.365 5.330 1.675 ;
        RECT  5.110 0.865 5.210 1.095 ;
        RECT  5.145 1.505 5.210 1.675 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  4.260 0.730 4.450 1.125 ;
        END
        AntennaGateArea 0.067 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.420 0.865 1.610 1.375 ;
        END
        AntennaGateArea 0.156 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.715 -0.210 6.160 0.210 ;
        RECT  5.545 -0.210 5.715 0.830 ;
        RECT  4.635 -0.210 5.545 0.210 ;
        RECT  4.465 -0.210 4.635 0.580 ;
        RECT  3.555 -0.210 4.465 0.210 ;
        RECT  3.385 -0.210 3.555 0.655 ;
        RECT  1.590 -0.210 3.385 0.210 ;
        RECT  1.330 -0.210 1.590 0.410 ;
        RECT  0.230 -0.210 1.330 0.210 ;
        RECT  0.070 -0.210 0.230 0.745 ;
        RECT  0.000 -0.210 0.070 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.740 2.310 6.160 2.730 ;
        RECT  5.480 2.130 5.740 2.730 ;
        RECT  4.640 2.310 5.480 2.730 ;
        RECT  4.380 2.220 4.640 2.730 ;
        RECT  3.725 2.310 4.380 2.730 ;
        RECT  3.465 2.220 3.725 2.730 ;
        RECT  1.880 2.310 3.465 2.730 ;
        RECT  1.620 2.220 1.880 2.730 ;
        RECT  0.230 2.310 1.620 2.730 ;
        RECT  0.070 1.520 0.230 2.730 ;
        RECT  0.000 2.310 0.070 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.760 1.015 5.810 1.275 ;
        RECT  5.640 1.015 5.760 2.010 ;
        RECT  4.990 1.890 5.640 2.010 ;
        RECT  4.870 0.425 4.990 2.100 ;
        RECT  4.810 0.425 4.870 0.895 ;
        RECT  4.830 1.430 4.870 2.100 ;
        RECT  3.335 1.980 4.830 2.100 ;
        RECT  4.690 1.010 4.750 1.270 ;
        RECT  4.570 1.010 4.690 1.860 ;
        RECT  0.950 1.740 4.570 1.860 ;
        RECT  4.140 0.420 4.255 0.590 ;
        RECT  4.140 1.260 4.230 1.600 ;
        RECT  4.110 0.420 4.140 1.600 ;
        RECT  4.020 0.420 4.110 1.380 ;
        RECT  3.580 1.210 4.020 1.380 ;
        RECT  2.250 1.500 3.960 1.620 ;
        RECT  3.770 0.440 3.890 1.015 ;
        RECT  2.250 0.895 3.770 1.015 ;
        RECT  2.430 1.260 3.580 1.380 ;
        RECT  3.165 1.980 3.335 2.150 ;
        RECT  2.770 1.980 3.030 2.135 ;
        RECT  0.590 1.980 2.770 2.100 ;
        RECT  2.480 0.505 2.740 0.690 ;
        RECT  1.060 0.570 2.480 0.690 ;
        RECT  2.130 0.895 2.250 1.620 ;
        RECT  1.190 1.500 2.130 1.620 ;
        RECT  1.070 1.215 1.190 1.620 ;
        RECT  1.025 1.215 1.070 1.335 ;
        RECT  0.940 0.570 1.060 0.920 ;
        RECT  0.855 1.085 1.025 1.335 ;
        RECT  0.830 1.500 0.950 1.860 ;
        RECT  0.660 0.330 0.940 0.450 ;
        RECT  0.710 0.800 0.940 0.920 ;
        RECT  0.710 1.500 0.830 1.620 ;
        RECT  0.590 0.800 0.710 1.620 ;
        RECT  0.540 0.330 0.660 0.640 ;
        RECT  0.470 1.780 0.590 2.100 ;
        RECT  0.470 0.520 0.540 0.640 ;
        RECT  0.350 0.520 0.470 1.900 ;
    END
END TLATNSRX2AD
MACRO TLATNSRX4AD
    CLASS CORE ;
    FOREIGN TLATNSRX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.280 0.980 0.510 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.970 0.910 5.110 1.030 ;
        RECT  4.850 0.910 4.970 1.380 ;
        RECT  3.850 1.260 4.850 1.380 ;
        RECT  3.700 1.145 3.850 1.380 ;
        RECT  3.580 0.900 3.700 1.380 ;
        RECT  2.740 0.900 3.580 1.020 ;
        RECT  2.480 0.900 2.740 1.070 ;
        END
        AntennaGateArea 0.269 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.330 0.375 8.500 1.590 ;
        RECT  8.190 1.005 8.330 1.590 ;
        END
        AntennaDiffArea 0.45 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.610 0.370 7.780 1.590 ;
        END
        AntennaDiffArea 0.422 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  6.350 0.785 6.650 1.105 ;
        END
        AntennaGateArea 0.1 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.180 1.140 3.440 1.330 ;
        RECT  2.085 1.210 3.180 1.330 ;
        RECT  1.690 1.130 2.085 1.330 ;
        END
        AntennaGateArea 0.296 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.870 -0.210 8.960 0.210 ;
        RECT  8.700 -0.210 8.870 0.860 ;
        RECT  8.135 -0.210 8.700 0.210 ;
        RECT  7.965 -0.210 8.135 0.860 ;
        RECT  7.395 -0.210 7.965 0.210 ;
        RECT  7.225 -0.210 7.395 0.560 ;
        RECT  6.640 -0.210 7.225 0.210 ;
        RECT  6.480 -0.210 6.640 0.660 ;
        RECT  5.595 -0.210 6.480 0.210 ;
        RECT  5.335 -0.210 5.595 0.310 ;
        RECT  3.240 -0.210 5.335 0.210 ;
        RECT  2.980 -0.210 3.240 0.300 ;
        RECT  1.655 -0.210 2.980 0.210 ;
        RECT  1.395 -0.210 1.655 0.300 ;
        RECT  0.840 -0.210 1.395 0.210 ;
        RECT  0.680 -0.210 0.840 0.610 ;
        RECT  0.000 -0.210 0.680 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.875 2.310 8.960 2.730 ;
        RECT  8.705 1.950 8.875 2.730 ;
        RECT  8.135 2.310 8.705 2.730 ;
        RECT  7.965 1.950 8.135 2.730 ;
        RECT  7.395 2.310 7.965 2.730 ;
        RECT  7.225 1.955 7.395 2.730 ;
        RECT  6.720 2.310 7.225 2.730 ;
        RECT  6.460 2.250 6.720 2.730 ;
        RECT  5.765 2.310 6.460 2.730 ;
        RECT  5.505 2.230 5.765 2.730 ;
        RECT  4.100 2.310 5.505 2.730 ;
        RECT  3.840 2.220 4.100 2.730 ;
        RECT  2.090 2.310 3.840 2.730 ;
        RECT  1.830 2.220 2.090 2.730 ;
        RECT  0.385 2.310 1.830 2.730 ;
        RECT  0.215 1.585 0.385 2.730 ;
        RECT  0.000 2.310 0.215 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.960 2.520 ;
        LAYER M1 ;
        RECT  8.670 1.040 8.790 1.830 ;
        RECT  7.445 1.710 8.670 1.830 ;
        RECT  7.325 0.680 7.445 1.830 ;
        RECT  7.005 0.680 7.325 0.800 ;
        RECT  7.070 1.710 7.325 1.830 ;
        RECT  6.980 1.085 7.200 1.255 ;
        RECT  7.030 1.645 7.070 1.830 ;
        RECT  6.885 1.645 7.030 2.100 ;
        RECT  6.835 0.625 7.005 0.800 ;
        RECT  6.770 1.085 6.980 1.410 ;
        RECT  5.220 1.980 6.885 2.100 ;
        RECT  6.700 1.255 6.770 1.410 ;
        RECT  6.580 1.255 6.700 1.860 ;
        RECT  1.140 1.740 6.580 1.860 ;
        RECT  6.230 1.260 6.335 1.620 ;
        RECT  6.230 0.430 6.285 0.650 ;
        RECT  6.215 0.430 6.230 1.620 ;
        RECT  6.110 0.430 6.215 1.380 ;
        RECT  5.115 0.430 6.110 0.550 ;
        RECT  5.600 0.930 6.110 1.190 ;
        RECT  5.370 1.500 6.065 1.620 ;
        RECT  5.370 0.670 5.990 0.790 ;
        RECT  5.250 0.670 5.370 1.620 ;
        RECT  4.700 0.670 5.250 0.790 ;
        RECT  3.220 1.500 5.250 1.620 ;
        RECT  4.995 0.400 5.115 0.550 ;
        RECT  4.840 1.980 5.100 2.190 ;
        RECT  4.460 0.400 4.995 0.520 ;
        RECT  3.220 1.980 4.840 2.100 ;
        RECT  4.580 0.640 4.700 0.900 ;
        RECT  4.340 0.400 4.460 0.780 ;
        RECT  4.200 0.660 4.340 0.780 ;
        RECT  1.125 0.420 4.220 0.540 ;
        RECT  4.080 0.660 4.200 1.140 ;
        RECT  1.870 0.660 4.080 0.780 ;
        RECT  2.960 1.450 3.220 1.620 ;
        RECT  2.940 1.980 3.220 2.190 ;
        RECT  1.380 1.500 2.960 1.620 ;
        RECT  0.810 1.980 2.940 2.100 ;
        RECT  1.750 0.660 1.870 0.930 ;
        RECT  1.260 1.040 1.380 1.620 ;
        RECT  1.170 1.040 1.260 1.320 ;
        RECT  1.050 1.440 1.140 1.860 ;
        RECT  1.050 0.420 1.125 0.900 ;
        RECT  1.005 0.420 1.050 1.860 ;
        RECT  0.930 0.780 1.005 1.860 ;
        RECT  0.690 0.735 0.810 2.100 ;
        RECT  0.385 0.735 0.690 0.855 ;
        RECT  0.575 1.585 0.690 2.100 ;
        RECT  0.215 0.345 0.385 0.855 ;
    END
END TLATNSRX4AD
MACRO TLATNSRXLAD
    CLASS CORE ;
    FOREIGN TLATNSRXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.855 0.230 1.375 ;
        END
        AntennaGateArea 0.053 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.910 1.935 1.330 ;
        END
        AntennaGateArea 0.091 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 0.670 5.530 1.800 ;
        RECT  5.335 0.670 5.390 0.840 ;
        RECT  5.335 1.630 5.390 1.800 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.830 0.490 4.970 1.750 ;
        RECT  4.620 0.490 4.830 0.610 ;
        RECT  4.680 1.490 4.830 1.750 ;
        END
        AntennaDiffArea 0.127 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.765 3.350 1.095 ;
        END
        AntennaGateArea 0.068 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.005 1.510 1.375 ;
        END
        AntennaGateArea 0.083 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.260 -0.210 5.600 0.210 ;
        RECT  5.000 -0.210 5.260 0.370 ;
        RECT  4.460 -0.210 5.000 0.210 ;
        RECT  4.200 -0.210 4.460 0.510 ;
        RECT  3.330 -0.210 4.200 0.210 ;
        RECT  3.070 -0.210 3.330 0.310 ;
        RECT  1.390 -0.210 3.070 0.210 ;
        RECT  1.130 -0.210 1.390 0.310 ;
        RECT  0.230 -0.210 1.130 0.210 ;
        RECT  0.070 -0.210 0.230 0.660 ;
        RECT  0.000 -0.210 0.070 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.170 2.310 5.600 2.730 ;
        RECT  4.910 2.215 5.170 2.730 ;
        RECT  4.220 2.310 4.910 2.730 ;
        RECT  3.960 2.220 4.220 2.730 ;
        RECT  3.235 2.310 3.960 2.730 ;
        RECT  2.975 1.975 3.235 2.730 ;
        RECT  1.680 2.310 2.975 2.730 ;
        RECT  1.420 2.215 1.680 2.730 ;
        RECT  0.360 2.310 1.420 2.730 ;
        RECT  0.100 2.210 0.360 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  5.210 0.990 5.270 1.250 ;
        RECT  5.090 0.990 5.210 2.095 ;
        RECT  4.560 1.975 5.090 2.095 ;
        RECT  4.560 0.760 4.680 1.020 ;
        RECT  4.440 0.760 4.560 2.095 ;
        RECT  3.835 1.975 4.440 2.095 ;
        RECT  4.200 1.110 4.320 1.855 ;
        RECT  0.825 1.735 4.200 1.855 ;
        RECT  3.960 0.445 4.080 1.615 ;
        RECT  3.880 0.445 3.960 0.705 ;
        RECT  2.190 1.495 3.960 1.615 ;
        RECT  3.665 0.830 3.840 1.090 ;
        RECT  3.575 1.975 3.835 2.190 ;
        RECT  3.530 0.435 3.665 1.365 ;
        RECT  3.495 0.435 3.530 0.605 ;
        RECT  3.470 1.085 3.530 1.365 ;
        RECT  2.570 1.245 3.470 1.365 ;
        RECT  2.310 1.200 2.570 1.365 ;
        RECT  2.190 0.900 2.560 1.020 ;
        RECT  2.210 0.590 2.350 0.710 ;
        RECT  2.090 0.455 2.210 0.710 ;
        RECT  1.940 1.975 2.200 2.190 ;
        RECT  2.070 0.900 2.190 1.615 ;
        RECT  1.120 0.455 2.090 0.575 ;
        RECT  1.070 1.495 2.070 1.615 ;
        RECT  0.555 1.975 1.940 2.095 ;
        RECT  1.000 0.455 1.120 0.830 ;
        RECT  0.950 0.960 1.070 1.615 ;
        RECT  0.710 0.710 1.000 0.830 ;
        RECT  0.830 0.960 0.950 1.220 ;
        RECT  0.750 0.330 0.870 0.590 ;
        RECT  0.710 1.380 0.825 1.855 ;
        RECT  0.470 0.470 0.750 0.590 ;
        RECT  0.705 0.710 0.710 1.855 ;
        RECT  0.590 0.710 0.705 1.550 ;
        RECT  0.470 1.730 0.555 2.095 ;
        RECT  0.435 0.470 0.470 2.095 ;
        RECT  0.350 0.470 0.435 1.900 ;
    END
END TLATNSRXLAD
MACRO TLATNTSCAX12AD
    CLASS CORE ;
    FOREIGN TLATNTSCAX12AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.955 0.960 2.170 1.375 ;
        END
        AntennaGateArea 0.109 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.940 0.380 11.310 2.130 ;
        RECT  8.460 0.380 10.940 0.540 ;
        RECT  10.840 1.125 10.940 2.130 ;
        RECT  10.025 1.440 10.840 1.820 ;
        RECT  9.855 1.440 10.025 2.130 ;
        RECT  8.775 1.440 9.855 1.820 ;
        RECT  8.605 1.440 8.775 2.170 ;
        END
        AntennaDiffArea 1.148 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.305 0.960 2.520 1.375 ;
        END
        AntennaGateArea 0.109 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.015 0.700 1.275 ;
        RECT  0.320 1.015 0.490 1.375 ;
        RECT  0.070 1.145 0.320 1.375 ;
        END
        AntennaGateArea 0.459 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.965 -0.210 11.480 0.210 ;
        RECT  10.705 -0.210 10.965 0.260 ;
        RECT  10.130 -0.210 10.705 0.210 ;
        RECT  9.610 -0.210 10.130 0.260 ;
        RECT  9.100 -0.210 9.610 0.210 ;
        RECT  8.840 -0.210 9.100 0.260 ;
        RECT  8.190 -0.210 8.840 0.210 ;
        RECT  7.670 -0.210 8.190 0.310 ;
        RECT  6.310 -0.210 7.670 0.210 ;
        RECT  6.050 -0.210 6.310 0.355 ;
        RECT  5.050 -0.210 6.050 0.210 ;
        RECT  4.790 -0.210 5.050 0.380 ;
        RECT  3.735 -0.210 4.790 0.210 ;
        RECT  3.475 -0.210 3.735 0.365 ;
        RECT  2.870 -0.210 3.475 0.210 ;
        RECT  2.610 -0.210 2.870 0.300 ;
        RECT  2.010 -0.210 2.610 0.210 ;
        RECT  1.750 -0.210 2.010 0.300 ;
        RECT  1.350 -0.210 1.750 0.210 ;
        RECT  1.190 -0.210 1.350 0.840 ;
        RECT  0.615 -0.210 1.190 0.210 ;
        RECT  0.445 -0.210 0.615 0.585 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  10.645 2.310 11.480 2.730 ;
        RECT  10.475 2.025 10.645 2.730 ;
        RECT  9.440 2.310 10.475 2.730 ;
        RECT  9.180 2.025 9.440 2.730 ;
        RECT  8.130 2.310 9.180 2.730 ;
        RECT  7.610 2.130 8.130 2.730 ;
        RECT  6.290 2.310 7.610 2.730 ;
        RECT  6.030 2.130 6.290 2.730 ;
        RECT  5.050 2.310 6.030 2.730 ;
        RECT  4.790 2.130 5.050 2.730 ;
        RECT  3.730 2.310 4.790 2.730 ;
        RECT  3.470 2.130 3.730 2.730 ;
        RECT  2.910 2.310 3.470 2.730 ;
        RECT  2.650 2.130 2.910 2.730 ;
        RECT  2.010 2.310 2.650 2.730 ;
        RECT  1.750 2.220 2.010 2.730 ;
        RECT  1.380 2.310 1.750 2.730 ;
        RECT  1.120 2.130 1.380 2.730 ;
        RECT  0.615 2.310 1.120 2.730 ;
        RECT  0.445 1.785 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 11.480 2.520 ;
        LAYER M1 ;
        RECT  10.200 0.870 10.820 0.990 ;
        RECT  10.080 0.660 10.200 1.260 ;
        RECT  8.340 0.660 10.080 0.780 ;
        RECT  8.680 1.140 10.080 1.260 ;
        RECT  8.290 0.900 9.690 1.020 ;
        RECT  8.220 0.435 8.340 0.780 ;
        RECT  8.170 0.900 8.290 2.010 ;
        RECT  7.310 0.435 8.220 0.555 ;
        RECT  7.090 1.890 8.170 2.010 ;
        RECT  7.890 0.680 8.010 1.520 ;
        RECT  7.800 1.400 7.890 1.520 ;
        RECT  7.550 1.400 7.800 1.620 ;
        RECT  7.650 0.990 7.770 1.250 ;
        RECT  7.310 0.990 7.650 1.110 ;
        RECT  7.430 1.360 7.550 1.620 ;
        RECT  7.190 0.435 7.310 1.755 ;
        RECT  4.160 0.510 7.190 0.630 ;
        RECT  4.160 1.635 7.190 1.755 ;
        RECT  6.830 1.890 7.090 2.190 ;
        RECT  6.950 0.750 7.070 1.470 ;
        RECT  4.040 0.750 6.950 0.870 ;
        RECT  4.290 1.350 6.950 1.470 ;
        RECT  4.040 1.890 6.830 2.010 ;
        RECT  4.040 1.050 6.810 1.170 ;
        RECT  3.920 0.490 4.040 0.870 ;
        RECT  3.920 1.050 4.040 2.010 ;
        RECT  3.280 0.490 3.920 0.610 ;
        RECT  0.980 1.890 3.920 2.010 ;
        RECT  3.645 0.730 3.800 1.475 ;
        RECT  3.030 0.730 3.645 0.850 ;
        RECT  3.280 1.355 3.645 1.475 ;
        RECT  2.890 1.060 3.365 1.230 ;
        RECT  3.160 0.420 3.280 0.610 ;
        RECT  3.130 1.355 3.280 1.750 ;
        RECT  1.670 0.420 3.160 0.540 ;
        RECT  3.020 1.630 3.130 1.750 ;
        RECT  2.770 0.660 2.890 1.770 ;
        RECT  2.130 0.660 2.770 0.780 ;
        RECT  2.425 1.600 2.770 1.770 ;
        RECT  1.670 1.590 1.740 1.710 ;
        RECT  1.550 0.420 1.670 1.710 ;
        RECT  1.480 1.590 1.550 1.710 ;
        RECT  0.980 1.020 1.430 1.280 ;
        RECT  0.975 1.020 0.980 2.010 ;
        RECT  0.830 0.400 0.975 2.010 ;
        RECT  0.255 0.750 0.830 0.870 ;
        RECT  0.255 1.545 0.830 1.665 ;
        RECT  0.085 0.375 0.255 0.870 ;
        RECT  0.085 1.545 0.255 2.080 ;
    END
END TLATNTSCAX12AD
MACRO TLATNTSCAX16AD
    CLASS CORE ;
    FOREIGN TLATNTSCAX16AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.035 2.855 1.375 ;
        END
        AntennaGateArea 0.144 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.645 0.385 12.990 1.970 ;
        RECT  12.520 0.385 12.645 2.115 ;
        RECT  8.910 0.385 12.520 0.715 ;
        RECT  12.475 1.125 12.520 2.115 ;
        RECT  12.090 1.125 12.475 1.970 ;
        RECT  11.410 1.470 12.090 1.970 ;
        RECT  11.240 1.470 11.410 2.160 ;
        RECT  10.190 1.470 11.240 1.970 ;
        RECT  10.020 1.470 10.190 2.180 ;
        RECT  8.970 1.470 10.020 1.970 ;
        RECT  8.800 1.470 8.970 2.160 ;
        END
        AntennaDiffArea 1.502 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.995 2.470 1.375 ;
        END
        AntennaGateArea 0.144 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.290 1.090 1.070 1.330 ;
        END
        AntennaGateArea 0.604 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.710 -0.210 13.160 0.210 ;
        RECT  12.450 -0.210 12.710 0.265 ;
        RECT  11.880 -0.210 12.450 0.210 ;
        RECT  11.360 -0.210 11.880 0.265 ;
        RECT  10.815 -0.210 11.360 0.210 ;
        RECT  10.295 -0.210 10.815 0.265 ;
        RECT  9.775 -0.210 10.295 0.210 ;
        RECT  9.255 -0.210 9.775 0.265 ;
        RECT  8.745 -0.210 9.255 0.210 ;
        RECT  8.485 -0.210 8.745 0.260 ;
        RECT  7.810 -0.210 8.485 0.210 ;
        RECT  7.550 -0.210 7.810 0.260 ;
        RECT  6.545 -0.210 7.550 0.210 ;
        RECT  6.285 -0.210 6.545 0.295 ;
        RECT  5.240 -0.210 6.285 0.210 ;
        RECT  4.980 -0.210 5.240 0.380 ;
        RECT  3.930 -0.210 4.980 0.210 ;
        RECT  3.670 -0.210 3.930 0.390 ;
        RECT  3.130 -0.210 3.670 0.210 ;
        RECT  2.870 -0.210 3.130 0.390 ;
        RECT  2.370 -0.210 2.870 0.210 ;
        RECT  2.110 -0.210 2.370 0.385 ;
        RECT  1.695 -0.210 2.110 0.210 ;
        RECT  1.525 -0.210 1.695 0.815 ;
        RECT  0.975 -0.210 1.525 0.210 ;
        RECT  0.805 -0.210 0.975 0.670 ;
        RECT  0.255 -0.210 0.805 0.210 ;
        RECT  0.085 -0.210 0.255 0.865 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  12.065 2.310 13.160 2.730 ;
        RECT  11.805 2.130 12.065 2.730 ;
        RECT  10.845 2.310 11.805 2.730 ;
        RECT  10.585 2.130 10.845 2.730 ;
        RECT  9.625 2.310 10.585 2.730 ;
        RECT  9.365 2.100 9.625 2.730 ;
        RECT  8.405 2.310 9.365 2.730 ;
        RECT  8.145 2.130 8.405 2.730 ;
        RECT  7.810 2.310 8.145 2.730 ;
        RECT  7.550 2.130 7.810 2.730 ;
        RECT  6.480 2.310 7.550 2.730 ;
        RECT  6.220 2.130 6.480 2.730 ;
        RECT  5.240 2.310 6.220 2.730 ;
        RECT  4.980 2.130 5.240 2.730 ;
        RECT  3.880 2.310 4.980 2.730 ;
        RECT  3.620 2.130 3.880 2.730 ;
        RECT  3.070 2.310 3.620 2.730 ;
        RECT  2.810 2.130 3.070 2.730 ;
        RECT  1.740 2.310 2.810 2.730 ;
        RECT  1.480 1.960 1.740 2.730 ;
        RECT  0.975 2.310 1.480 2.730 ;
        RECT  0.805 1.795 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.565 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 13.160 2.520 ;
        LAYER M1 ;
        RECT  8.790 0.885 12.390 1.005 ;
        RECT  8.485 1.135 11.945 1.255 ;
        RECT  8.670 0.380 8.790 1.005 ;
        RECT  7.525 0.380 8.670 0.500 ;
        RECT  8.365 1.040 8.485 2.010 ;
        RECT  7.280 1.890 8.365 2.010 ;
        RECT  8.100 0.680 8.220 1.520 ;
        RECT  8.010 1.400 8.100 1.520 ;
        RECT  7.645 1.400 8.010 1.660 ;
        RECT  7.860 0.990 7.980 1.250 ;
        RECT  7.525 0.990 7.860 1.110 ;
        RECT  7.405 0.380 7.525 1.755 ;
        RECT  4.300 0.510 7.405 0.630 ;
        RECT  4.350 1.635 7.405 1.755 ;
        RECT  7.165 0.790 7.285 1.470 ;
        RECT  7.020 1.890 7.280 2.190 ;
        RECT  4.175 0.790 7.165 0.910 ;
        RECT  4.470 1.350 7.165 1.470 ;
        RECT  6.785 1.030 7.045 1.190 ;
        RECT  4.190 1.890 7.020 2.010 ;
        RECT  4.190 1.070 6.785 1.190 ;
        RECT  4.070 1.070 4.190 2.010 ;
        RECT  4.055 0.510 4.175 0.910 ;
        RECT  1.980 1.890 4.070 2.010 ;
        RECT  2.030 0.510 4.055 0.630 ;
        RECT  3.660 1.040 3.950 1.300 ;
        RECT  3.540 0.750 3.660 1.770 ;
        RECT  3.230 0.750 3.540 0.870 ;
        RECT  3.260 1.510 3.540 1.770 ;
        RECT  3.110 1.040 3.230 1.300 ;
        RECT  2.990 0.750 3.110 1.770 ;
        RECT  2.490 0.750 2.990 0.870 ;
        RECT  2.180 1.650 2.990 1.770 ;
        RECT  1.910 0.510 2.030 1.600 ;
        RECT  1.860 1.720 1.980 2.010 ;
        RECT  1.310 1.720 1.860 1.840 ;
        RECT  1.310 1.020 1.790 1.280 ;
        RECT  1.190 0.390 1.310 2.040 ;
        RECT  0.590 0.790 1.190 0.910 ;
        RECT  0.590 1.520 1.190 1.640 ;
        RECT  0.470 0.390 0.590 0.910 ;
        RECT  0.470 1.520 0.590 2.040 ;
    END
END TLATNTSCAX16AD
MACRO TLATNTSCAX20AD
    CLASS CORE ;
    FOREIGN TLATNTSCAX20AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.340 1.040 3.460 1.375 ;
        RECT  3.150 1.110 3.340 1.375 ;
        END
        AntennaGateArea 0.158 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.500 0.415 16.100 2.010 ;
        RECT  10.630 0.415 15.500 0.715 ;
        RECT  15.170 1.125 15.500 2.010 ;
        RECT  14.515 1.430 15.170 2.010 ;
        RECT  14.345 1.430 14.515 2.145 ;
        RECT  13.235 1.430 14.345 2.010 ;
        RECT  13.065 1.430 13.235 2.140 ;
        RECT  11.975 1.430 13.065 2.010 ;
        RECT  11.805 1.430 11.975 2.135 ;
        RECT  10.745 1.430 11.805 2.010 ;
        RECT  10.575 1.430 10.745 2.135 ;
        END
        AntennaDiffArea 1.808 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.730 1.040 2.790 1.375 ;
        RECT  2.590 0.865 2.730 1.375 ;
        END
        AntennaGateArea 0.158 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.300 1.130 1.340 1.330 ;
        END
        AntennaGateArea 0.755 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.620 -0.210 16.240 0.210 ;
        RECT  15.360 -0.210 15.620 0.280 ;
        RECT  14.675 -0.210 15.360 0.210 ;
        RECT  14.415 -0.210 14.675 0.295 ;
        RECT  13.670 -0.210 14.415 0.210 ;
        RECT  13.150 -0.210 13.670 0.295 ;
        RECT  12.510 -0.210 13.150 0.210 ;
        RECT  11.990 -0.210 12.510 0.290 ;
        RECT  11.310 -0.210 11.990 0.210 ;
        RECT  11.050 -0.210 11.310 0.290 ;
        RECT  10.440 -0.210 11.050 0.210 ;
        RECT  10.180 -0.210 10.440 0.300 ;
        RECT  9.720 -0.210 10.180 0.210 ;
        RECT  9.460 -0.210 9.720 0.265 ;
        RECT  8.885 -0.210 9.460 0.210 ;
        RECT  8.625 -0.210 8.885 0.300 ;
        RECT  7.580 -0.210 8.625 0.210 ;
        RECT  7.320 -0.210 7.580 0.425 ;
        RECT  6.320 -0.210 7.320 0.210 ;
        RECT  6.060 -0.210 6.320 0.425 ;
        RECT  5.060 -0.210 6.060 0.210 ;
        RECT  4.800 -0.210 5.060 0.230 ;
        RECT  4.430 -0.210 4.800 0.210 ;
        RECT  4.170 -0.210 4.430 0.300 ;
        RECT  3.670 -0.210 4.170 0.210 ;
        RECT  3.410 -0.210 3.670 0.300 ;
        RECT  2.810 -0.210 3.410 0.210 ;
        RECT  2.550 -0.210 2.810 0.300 ;
        RECT  2.120 -0.210 2.550 0.210 ;
        RECT  1.860 -0.210 2.120 0.270 ;
        RECT  1.380 -0.210 1.860 0.210 ;
        RECT  1.120 -0.210 1.380 0.650 ;
        RECT  0.660 -0.210 1.120 0.210 ;
        RECT  0.400 -0.210 0.660 0.650 ;
        RECT  0.000 -0.210 0.400 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  15.180 2.310 16.240 2.730 ;
        RECT  14.920 2.130 15.180 2.730 ;
        RECT  13.920 2.310 14.920 2.730 ;
        RECT  13.660 2.130 13.920 2.730 ;
        RECT  12.650 2.310 13.660 2.730 ;
        RECT  12.390 2.130 12.650 2.730 ;
        RECT  11.400 2.310 12.390 2.730 ;
        RECT  11.140 2.130 11.400 2.730 ;
        RECT  10.100 2.310 11.140 2.730 ;
        RECT  9.580 2.130 10.100 2.730 ;
        RECT  8.820 2.310 9.580 2.730 ;
        RECT  8.560 2.130 8.820 2.730 ;
        RECT  7.600 2.310 8.560 2.730 ;
        RECT  7.340 2.130 7.600 2.730 ;
        RECT  6.340 2.310 7.340 2.730 ;
        RECT  6.080 2.130 6.340 2.730 ;
        RECT  5.080 2.310 6.080 2.730 ;
        RECT  4.820 2.130 5.080 2.730 ;
        RECT  4.430 2.310 4.820 2.730 ;
        RECT  4.170 2.190 4.430 2.730 ;
        RECT  3.670 2.310 4.170 2.730 ;
        RECT  3.410 2.130 3.670 2.730 ;
        RECT  2.700 2.310 3.410 2.730 ;
        RECT  2.440 2.220 2.700 2.730 ;
        RECT  2.120 2.310 2.440 2.730 ;
        RECT  1.860 2.220 2.120 2.730 ;
        RECT  1.335 2.310 1.860 2.730 ;
        RECT  1.165 1.795 1.335 2.730 ;
        RECT  0.615 2.310 1.165 2.730 ;
        RECT  0.445 1.795 0.615 2.730 ;
        RECT  0.000 2.310 0.445 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 16.240 2.520 ;
        LAYER M1 ;
        RECT  10.510 0.885 15.375 1.005 ;
        RECT  10.260 1.140 15.050 1.260 ;
        RECT  10.390 0.450 10.510 1.005 ;
        RECT  9.180 0.450 10.390 0.570 ;
        RECT  10.140 1.040 10.260 2.010 ;
        RECT  9.215 1.890 10.140 2.010 ;
        RECT  10.020 0.690 10.100 0.810 ;
        RECT  9.900 0.690 10.020 1.460 ;
        RECT  9.840 0.690 9.900 0.810 ;
        RECT  9.760 1.340 9.900 1.460 ;
        RECT  9.660 0.940 9.780 1.200 ;
        RECT  9.640 1.340 9.760 1.620 ;
        RECT  9.180 1.010 9.660 1.130 ;
        RECT  9.495 1.340 9.640 1.460 ;
        RECT  9.375 1.280 9.495 1.540 ;
        RECT  8.955 1.890 9.215 2.050 ;
        RECT  9.060 0.450 9.180 1.770 ;
        RECT  8.940 0.545 9.060 0.840 ;
        RECT  5.470 1.650 9.060 1.770 ;
        RECT  5.200 1.890 8.955 2.010 ;
        RECT  5.430 0.545 8.940 0.665 ;
        RECT  8.780 0.995 8.940 1.255 ;
        RECT  8.660 0.785 8.780 1.470 ;
        RECT  5.250 0.785 8.660 0.905 ;
        RECT  5.580 1.350 8.660 1.470 ;
        RECT  5.400 1.070 8.385 1.190 ;
        RECT  5.280 1.070 5.400 1.540 ;
        RECT  5.200 1.420 5.280 1.540 ;
        RECT  5.130 0.420 5.250 0.905 ;
        RECT  5.080 1.420 5.200 2.010 ;
        RECT  4.740 1.040 5.160 1.300 ;
        RECT  2.460 0.420 5.130 0.540 ;
        RECT  1.670 1.890 5.080 2.010 ;
        RECT  4.740 0.760 4.810 0.880 ;
        RECT  4.620 0.760 4.740 1.770 ;
        RECT  3.785 0.760 4.620 0.880 ;
        RECT  3.980 1.650 4.620 1.770 ;
        RECT  3.720 1.050 4.380 1.310 ;
        RECT  3.860 1.510 3.980 1.770 ;
        RECT  3.580 1.050 3.720 1.770 ;
        RECT  3.030 1.650 3.580 1.770 ;
        RECT  3.030 0.660 3.290 0.780 ;
        RECT  2.910 0.660 3.030 1.770 ;
        RECT  2.780 1.650 2.910 1.770 ;
        RECT  2.340 0.420 2.460 1.730 ;
        RECT  2.220 0.620 2.340 0.880 ;
        RECT  2.220 1.470 2.340 1.730 ;
        RECT  1.670 1.070 2.220 1.190 ;
        RECT  1.550 0.370 1.670 2.010 ;
        RECT  0.950 0.770 1.550 0.890 ;
        RECT  0.975 1.520 1.550 1.640 ;
        RECT  0.805 1.520 0.975 1.995 ;
        RECT  0.830 0.370 0.950 0.890 ;
        RECT  0.230 0.770 0.830 0.890 ;
        RECT  0.255 1.520 0.805 1.640 ;
        RECT  0.085 1.520 0.255 1.995 ;
        RECT  0.110 0.370 0.230 0.890 ;
    END
END TLATNTSCAX20AD
MACRO TLATNTSCAX2AD
    CLASS CORE ;
    FOREIGN TLATNTSCAX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.400 1.090 1.610 1.375 ;
        RECT  1.280 0.950 1.400 1.375 ;
        END
        AntennaGateArea 0.055 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.770 1.425 4.920 2.030 ;
        RECT  4.700 1.425 4.770 1.655 ;
        RECT  4.550 0.760 4.700 1.655 ;
        RECT  4.440 0.760 4.550 0.880 ;
        END
        AntennaDiffArea 0.276 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.730 0.965 1.890 1.375 ;
        END
        AntennaGateArea 0.055 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.020 0.235 1.375 ;
        END
        AntennaGateArea 0.114 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.930 -0.210 5.040 0.210 ;
        RECT  4.670 -0.210 4.930 0.395 ;
        RECT  4.410 -0.210 4.670 0.210 ;
        RECT  4.150 -0.210 4.410 0.395 ;
        RECT  3.865 -0.210 4.150 0.210 ;
        RECT  3.605 -0.210 3.865 0.390 ;
        RECT  2.405 -0.210 3.605 0.210 ;
        RECT  1.885 -0.210 2.405 0.330 ;
        RECT  1.095 -0.210 1.885 0.210 ;
        RECT  0.475 -0.210 1.095 0.300 ;
        RECT  0.000 -0.210 0.475 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.295 2.310 5.040 2.730 ;
        RECT  3.775 2.130 4.295 2.730 ;
        RECT  2.495 2.310 3.775 2.730 ;
        RECT  2.235 2.220 2.495 2.730 ;
        RECT  1.235 2.310 2.235 2.730 ;
        RECT  0.975 2.050 1.235 2.730 ;
        RECT  0.680 2.310 0.975 2.730 ;
        RECT  0.420 2.030 0.680 2.730 ;
        RECT  0.000 2.310 0.420 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.040 2.520 ;
        LAYER M1 ;
        RECT  4.830 0.520 4.950 1.280 ;
        RECT  3.485 0.520 4.830 0.640 ;
        RECT  4.400 1.020 4.430 1.280 ;
        RECT  4.280 1.020 4.400 2.010 ;
        RECT  3.540 1.890 4.280 2.010 ;
        RECT  4.040 0.760 4.160 1.620 ;
        RECT  3.810 0.760 4.040 0.880 ;
        RECT  3.790 1.400 4.040 1.620 ;
        RECT  3.485 1.060 3.920 1.180 ;
        RECT  3.470 1.500 3.790 1.620 ;
        RECT  3.420 1.890 3.540 2.140 ;
        RECT  3.365 0.380 3.485 1.340 ;
        RECT  3.395 2.020 3.420 2.140 ;
        RECT  3.135 2.020 3.395 2.190 ;
        RECT  3.085 0.380 3.365 0.500 ;
        RECT  3.090 1.220 3.365 1.340 ;
        RECT  3.120 0.620 3.240 1.100 ;
        RECT  3.090 1.780 3.230 1.900 ;
        RECT  2.840 2.020 3.135 2.140 ;
        RECT  2.715 0.620 3.120 0.740 ;
        RECT  2.970 1.220 3.090 1.900 ;
        RECT  2.915 0.330 3.085 0.500 ;
        RECT  2.840 0.940 2.980 1.060 ;
        RECT  2.720 0.940 2.840 2.140 ;
        RECT  1.560 1.980 2.720 2.100 ;
        RECT  2.595 0.470 2.715 0.740 ;
        RECT  2.480 0.980 2.600 1.860 ;
        RECT  0.910 0.470 2.595 0.590 ;
        RECT  2.175 0.980 2.480 1.100 ;
        RECT  1.955 1.740 2.480 1.860 ;
        RECT  2.145 1.260 2.295 1.620 ;
        RECT  2.055 0.710 2.175 1.100 ;
        RECT  1.805 1.500 2.145 1.620 ;
        RECT  1.915 0.710 2.055 0.830 ;
        RECT  1.685 1.500 1.805 1.760 ;
        RECT  1.160 1.500 1.685 1.620 ;
        RECT  1.160 0.710 1.640 0.830 ;
        RECT  1.440 1.790 1.560 2.100 ;
        RECT  0.490 1.790 1.440 1.910 ;
        RECT  1.040 0.710 1.160 1.620 ;
        RECT  0.790 0.470 0.910 1.600 ;
        RECT  0.725 1.430 0.790 1.600 ;
        RECT  0.370 0.780 0.490 1.910 ;
        RECT  0.255 0.780 0.370 0.900 ;
        RECT  0.230 1.530 0.370 1.910 ;
        RECT  0.085 0.455 0.255 0.900 ;
        RECT  0.110 1.530 0.230 2.050 ;
    END
END TLATNTSCAX2AD
MACRO TLATNTSCAX3AD
    CLASS CORE ;
    FOREIGN TLATNTSCAX3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.140 0.710 1.330 1.095 ;
        END
        AntennaGateArea 0.055 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.750 1.425 4.970 1.810 ;
        RECT  4.750 0.750 4.820 0.870 ;
        RECT  4.630 0.750 4.750 1.810 ;
        RECT  4.560 0.750 4.630 0.870 ;
        END
        AntennaDiffArea 0.278 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 1.290 1.655 1.610 ;
        END
        AntennaGateArea 0.055 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.115 0.235 1.375 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.137 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.300 -0.210 5.600 0.210 ;
        RECT  5.180 -0.210 5.300 0.905 ;
        RECT  4.375 -0.210 5.180 0.210 ;
        RECT  3.685 -0.210 4.375 0.300 ;
        RECT  2.390 -0.210 3.685 0.210 ;
        RECT  1.870 -0.210 2.390 0.300 ;
        RECT  1.225 -0.210 1.870 0.210 ;
        RECT  0.445 -0.210 1.225 0.300 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.520 2.310 5.600 2.730 ;
        RECT  5.360 1.685 5.520 2.730 ;
        RECT  4.255 2.310 5.360 2.730 ;
        RECT  3.735 2.220 4.255 2.730 ;
        RECT  2.470 2.310 3.735 2.730 ;
        RECT  2.210 2.220 2.470 2.730 ;
        RECT  1.120 2.310 2.210 2.730 ;
        RECT  0.600 2.170 1.120 2.730 ;
        RECT  0.000 2.310 0.600 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  5.210 1.250 5.330 1.560 ;
        RECT  5.090 1.435 5.210 2.050 ;
        RECT  4.510 1.930 5.090 2.050 ;
        RECT  4.940 0.470 5.060 1.285 ;
        RECT  3.565 0.470 4.940 0.590 ;
        RECT  4.900 0.990 4.940 1.285 ;
        RECT  4.390 1.010 4.510 2.050 ;
        RECT  3.425 1.930 4.390 2.050 ;
        RECT  4.150 0.760 4.270 1.630 ;
        RECT  3.810 0.760 4.150 0.880 ;
        RECT  3.920 1.510 4.150 1.630 ;
        RECT  3.910 1.055 4.030 1.315 ;
        RECT  3.775 1.510 3.920 1.770 ;
        RECT  3.565 1.055 3.910 1.180 ;
        RECT  3.655 1.330 3.775 1.770 ;
        RECT  3.485 1.330 3.655 1.470 ;
        RECT  3.445 0.420 3.565 1.180 ;
        RECT  2.925 0.420 3.445 0.540 ;
        RECT  3.350 1.055 3.445 1.180 ;
        RECT  3.390 1.930 3.425 2.140 ;
        RECT  3.270 1.605 3.390 2.140 ;
        RECT  3.230 1.055 3.350 1.400 ;
        RECT  3.150 0.660 3.325 0.920 ;
        RECT  2.790 2.020 3.270 2.140 ;
        RECT  3.115 1.280 3.230 1.400 ;
        RECT  2.700 0.660 3.150 0.780 ;
        RECT  2.995 1.280 3.115 1.875 ;
        RECT  2.860 0.900 2.960 1.160 ;
        RECT  2.790 0.900 2.860 1.560 ;
        RECT  2.740 0.900 2.790 2.140 ;
        RECT  2.670 1.440 2.740 2.140 ;
        RECT  2.580 0.470 2.700 0.780 ;
        RECT  1.470 1.980 2.670 2.100 ;
        RECT  2.405 1.020 2.620 1.280 ;
        RECT  0.920 0.470 2.580 0.590 ;
        RECT  2.285 0.810 2.405 1.560 ;
        RECT  1.960 0.810 2.285 0.930 ;
        RECT  2.160 1.440 2.285 1.560 ;
        RECT  1.895 1.050 2.165 1.310 ;
        RECT  2.040 1.440 2.160 1.700 ;
        RECT  1.775 1.050 1.895 1.850 ;
        RECT  1.570 1.050 1.775 1.170 ;
        RECT  1.610 1.730 1.775 1.850 ;
        RECT  1.450 0.710 1.570 1.170 ;
        RECT  1.350 1.930 1.470 2.100 ;
        RECT  0.490 1.930 1.350 2.050 ;
        RECT  0.800 0.470 0.920 1.630 ;
        RECT  0.735 1.460 0.800 1.630 ;
        RECT  0.490 1.000 0.680 1.260 ;
        RECT  0.370 0.625 0.490 2.050 ;
        RECT  0.230 0.625 0.370 0.745 ;
        RECT  0.230 1.610 0.370 1.730 ;
        RECT  0.110 0.485 0.230 0.745 ;
        RECT  0.110 1.610 0.230 2.130 ;
    END
END TLATNTSCAX3AD
MACRO TLATNTSCAX4AD
    CLASS CORE ;
    FOREIGN TLATNTSCAX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.440 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.190 0.790 1.330 1.350 ;
        END
        AntennaGateArea 0.065 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.720 1.285 5.810 1.795 ;
        RECT  5.670 1.285 5.720 1.860 ;
        RECT  5.600 0.620 5.670 1.860 ;
        RECT  5.550 0.620 5.600 1.455 ;
        RECT  5.410 0.620 5.550 0.740 ;
        END
        AntennaDiffArea 0.428 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.470 1.670 1.610 ;
        RECT  1.520 1.265 1.640 1.610 ;
        RECT  1.145 1.470 1.520 1.610 ;
        END
        AntennaGateArea 0.065 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.240 1.010 0.335 1.270 ;
        RECT  0.070 0.865 0.240 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.150 -0.210 6.440 0.210 ;
        RECT  6.030 -0.210 6.150 0.630 ;
        RECT  5.290 -0.210 6.030 0.210 ;
        RECT  5.030 -0.210 5.290 0.245 ;
        RECT  4.660 -0.210 5.030 0.210 ;
        RECT  4.400 -0.210 4.660 0.260 ;
        RECT  3.770 -0.210 4.400 0.210 ;
        RECT  3.510 -0.210 3.770 0.260 ;
        RECT  2.410 -0.210 3.510 0.210 ;
        RECT  1.890 -0.210 2.410 0.245 ;
        RECT  1.120 -0.210 1.890 0.210 ;
        RECT  0.600 -0.210 1.120 0.300 ;
        RECT  0.000 -0.210 0.600 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.370 2.310 6.440 2.730 ;
        RECT  6.210 1.565 6.370 2.730 ;
        RECT  5.060 2.310 6.210 2.730 ;
        RECT  4.540 2.245 5.060 2.730 ;
        RECT  3.770 2.310 4.540 2.730 ;
        RECT  3.510 2.270 3.770 2.730 ;
        RECT  2.510 2.310 3.510 2.730 ;
        RECT  2.250 2.270 2.510 2.730 ;
        RECT  1.080 2.310 2.250 2.730 ;
        RECT  0.560 2.130 1.080 2.730 ;
        RECT  0.000 2.310 0.560 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.440 2.520 ;
        LAYER M1 ;
        RECT  6.165 1.070 6.285 1.335 ;
        RECT  6.090 1.215 6.165 1.335 ;
        RECT  5.970 1.215 6.090 2.110 ;
        RECT  5.160 1.980 5.970 2.110 ;
        RECT  5.790 0.380 5.910 1.090 ;
        RECT  5.210 0.380 5.790 0.500 ;
        RECT  5.160 1.140 5.300 1.260 ;
        RECT  5.090 0.380 5.210 0.980 ;
        RECT  5.040 1.140 5.160 2.110 ;
        RECT  4.300 0.380 5.090 0.500 ;
        RECT  4.900 0.860 5.090 0.980 ;
        RECT  4.140 1.990 5.040 2.110 ;
        RECT  4.600 0.620 4.910 0.740 ;
        RECT  4.780 0.860 4.900 1.215 ;
        RECT  4.600 1.400 4.820 1.520 ;
        RECT  4.480 0.620 4.600 1.520 ;
        RECT  4.170 0.380 4.300 1.805 ;
        RECT  3.095 0.560 4.170 0.680 ;
        RECT  4.020 1.685 4.170 1.805 ;
        RECT  3.880 1.990 4.140 2.165 ;
        RECT  3.760 1.685 4.020 1.870 ;
        RECT  2.740 1.990 3.880 2.110 ;
        RECT  3.650 0.800 3.770 1.490 ;
        RECT  3.070 1.685 3.760 1.805 ;
        RECT  2.805 0.800 3.650 0.920 ;
        RECT  3.000 1.370 3.650 1.490 ;
        RECT  2.925 0.510 3.095 0.680 ;
        RECT  2.950 1.610 3.070 1.870 ;
        RECT  2.855 1.060 3.020 1.180 ;
        RECT  2.740 1.060 2.855 1.535 ;
        RECT  2.685 0.470 2.805 0.920 ;
        RECT  2.735 1.060 2.740 2.110 ;
        RECT  2.620 1.415 2.735 2.110 ;
        RECT  0.920 0.470 2.685 0.590 ;
        RECT  1.475 1.990 2.620 2.110 ;
        RECT  2.500 1.035 2.610 1.295 ;
        RECT  2.380 0.825 2.500 1.655 ;
        RECT  2.175 0.825 2.380 0.945 ;
        RECT  2.150 1.535 2.380 1.655 ;
        RECT  1.910 1.065 2.260 1.325 ;
        RECT  2.005 0.710 2.175 0.945 ;
        RECT  2.030 1.535 2.150 1.795 ;
        RECT  1.885 1.065 1.910 1.860 ;
        RECT  1.790 0.850 1.885 1.860 ;
        RECT  1.765 0.850 1.790 1.185 ;
        RECT  1.610 1.740 1.790 1.860 ;
        RECT  1.570 0.850 1.765 0.970 ;
        RECT  1.450 0.710 1.570 0.970 ;
        RECT  1.355 1.780 1.475 2.110 ;
        RECT  0.585 1.780 1.355 1.900 ;
        RECT  0.800 0.470 0.920 1.650 ;
        RECT  0.715 1.480 0.800 1.650 ;
        RECT  0.585 1.000 0.680 1.260 ;
        RECT  0.465 0.625 0.585 1.900 ;
        RECT  0.255 0.625 0.465 0.745 ;
        RECT  0.255 1.750 0.465 1.900 ;
        RECT  0.085 0.465 0.255 0.745 ;
        RECT  0.085 1.575 0.255 2.005 ;
    END
END TLATNTSCAX4AD
MACRO TLATNTSCAX6AD
    CLASS CORE ;
    FOREIGN TLATNTSCAX6AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 0.960 1.750 1.220 ;
        RECT  1.470 0.865 1.610 1.375 ;
        END
        AntennaGateArea 0.058 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.125 0.380 8.245 1.675 ;
        RECT  8.065 0.380 8.125 2.175 ;
        RECT  6.545 0.380 8.065 0.540 ;
        RECT  7.925 1.430 8.065 2.175 ;
        RECT  6.865 1.430 7.925 1.610 ;
        RECT  6.665 1.430 6.865 2.175 ;
        END
        AntennaDiffArea 0.668 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.945 1.200 2.060 1.460 ;
        RECT  1.940 1.200 1.945 1.655 ;
        RECT  1.745 1.340 1.940 1.655 ;
        END
        AntennaGateArea 0.058 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.015 0.325 1.275 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.24 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.945 -0.210 8.400 0.210 ;
        RECT  7.685 -0.210 7.945 0.260 ;
        RECT  7.185 -0.210 7.685 0.210 ;
        RECT  6.925 -0.210 7.185 0.260 ;
        RECT  6.275 -0.210 6.925 0.210 ;
        RECT  5.755 -0.210 6.275 0.310 ;
        RECT  4.390 -0.210 5.755 0.210 ;
        RECT  4.130 -0.210 4.390 0.380 ;
        RECT  3.130 -0.210 4.130 0.210 ;
        RECT  2.870 -0.210 3.130 0.390 ;
        RECT  2.400 -0.210 2.870 0.210 ;
        RECT  2.140 -0.210 2.400 0.300 ;
        RECT  1.690 -0.210 2.140 0.210 ;
        RECT  1.430 -0.210 1.690 0.300 ;
        RECT  0.970 -0.210 1.430 0.210 ;
        RECT  0.810 -0.210 0.970 0.860 ;
        RECT  0.255 -0.210 0.810 0.210 ;
        RECT  0.085 -0.210 0.255 0.745 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.480 2.310 8.400 2.730 ;
        RECT  7.310 1.845 7.480 2.730 ;
        RECT  6.215 2.310 7.310 2.730 ;
        RECT  5.695 2.130 6.215 2.730 ;
        RECT  4.390 2.310 5.695 2.730 ;
        RECT  4.130 2.115 4.390 2.730 ;
        RECT  3.070 2.310 4.130 2.730 ;
        RECT  2.810 2.190 3.070 2.730 ;
        RECT  1.610 2.310 2.810 2.730 ;
        RECT  0.830 2.220 1.610 2.730 ;
        RECT  0.250 2.310 0.830 2.730 ;
        RECT  0.090 1.550 0.250 2.730 ;
        RECT  0.000 2.310 0.090 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.400 2.520 ;
        LAYER M1 ;
        RECT  7.825 0.660 7.945 1.260 ;
        RECT  6.425 0.660 7.825 0.780 ;
        RECT  6.765 1.140 7.825 1.260 ;
        RECT  6.375 0.900 7.685 1.020 ;
        RECT  6.305 0.435 6.425 0.780 ;
        RECT  6.255 0.900 6.375 1.995 ;
        RECT  5.385 0.435 6.305 0.555 ;
        RECT  5.325 1.875 6.255 1.995 ;
        RECT  5.975 0.690 6.095 1.520 ;
        RECT  5.885 1.400 5.975 1.520 ;
        RECT  5.625 1.400 5.885 1.655 ;
        RECT  5.735 1.000 5.855 1.260 ;
        RECT  5.385 1.075 5.735 1.195 ;
        RECT  5.505 1.355 5.625 1.655 ;
        RECT  5.265 0.435 5.385 1.755 ;
        RECT  5.065 1.875 5.325 2.190 ;
        RECT  3.500 0.510 5.265 0.630 ;
        RECT  3.500 1.635 5.265 1.755 ;
        RECT  5.020 0.750 5.140 1.470 ;
        RECT  3.380 1.875 5.065 1.995 ;
        RECT  3.375 0.750 5.020 0.870 ;
        RECT  3.630 1.350 5.020 1.470 ;
        RECT  3.380 1.050 4.900 1.170 ;
        RECT  3.260 1.050 3.380 2.050 ;
        RECT  3.255 0.510 3.375 0.870 ;
        RECT  0.590 1.930 3.260 2.050 ;
        RECT  2.705 0.510 3.255 0.630 ;
        RECT  3.065 1.215 3.140 1.475 ;
        RECT  2.945 0.750 3.065 1.475 ;
        RECT  2.490 0.750 2.945 0.870 ;
        RECT  2.550 1.355 2.945 1.475 ;
        RECT  2.310 1.060 2.825 1.230 ;
        RECT  2.585 0.420 2.705 0.630 ;
        RECT  1.310 0.420 2.585 0.540 ;
        RECT  2.430 1.355 2.550 1.765 ;
        RECT  2.190 0.660 2.310 1.810 ;
        RECT  1.810 0.660 2.190 0.780 ;
        RECT  2.065 1.640 2.190 1.810 ;
        RECT  1.190 0.420 1.310 1.725 ;
        RECT  1.115 1.555 1.190 1.725 ;
        RECT  0.590 1.020 1.070 1.280 ;
        RECT  0.470 0.400 0.590 2.050 ;
    END
END TLATNTSCAX6AD
MACRO TLATNTSCAX8AD
    CLASS CORE ;
    FOREIGN TLATNTSCAX8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.610 0.960 1.750 1.220 ;
        RECT  1.470 0.865 1.610 1.375 ;
        END
        AntennaGateArea 0.076 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.060 0.380 9.310 1.795 ;
        RECT  7.240 0.380 9.060 0.540 ;
        RECT  8.885 1.285 9.060 1.795 ;
        RECT  8.820 1.430 8.885 1.795 ;
        RECT  8.620 1.430 8.820 2.175 ;
        RECT  7.560 1.430 8.620 1.680 ;
        RECT  7.360 1.430 7.560 2.175 ;
        END
        AntennaDiffArea 0.768 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.945 1.200 2.060 1.460 ;
        RECT  1.940 1.200 1.945 1.655 ;
        RECT  1.745 1.340 1.940 1.655 ;
        END
        AntennaGateArea 0.076 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.015 0.325 1.275 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.312 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.640 -0.210 9.520 0.210 ;
        RECT  8.380 -0.210 8.640 0.260 ;
        RECT  7.880 -0.210 8.380 0.210 ;
        RECT  7.620 -0.210 7.880 0.260 ;
        RECT  6.970 -0.210 7.620 0.210 ;
        RECT  6.450 -0.210 6.970 0.310 ;
        RECT  5.660 -0.210 6.450 0.210 ;
        RECT  5.400 -0.210 5.660 0.355 ;
        RECT  4.390 -0.210 5.400 0.210 ;
        RECT  4.130 -0.210 4.390 0.380 ;
        RECT  3.130 -0.210 4.130 0.210 ;
        RECT  2.870 -0.210 3.130 0.390 ;
        RECT  2.400 -0.210 2.870 0.210 ;
        RECT  2.140 -0.210 2.400 0.300 ;
        RECT  1.690 -0.210 2.140 0.210 ;
        RECT  1.430 -0.210 1.690 0.300 ;
        RECT  0.970 -0.210 1.430 0.210 ;
        RECT  0.810 -0.210 0.970 0.840 ;
        RECT  0.255 -0.210 0.810 0.210 ;
        RECT  0.085 -0.210 0.255 0.745 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  9.425 2.310 9.520 2.730 ;
        RECT  9.255 2.025 9.425 2.730 ;
        RECT  8.220 2.310 9.255 2.730 ;
        RECT  7.960 1.870 8.220 2.730 ;
        RECT  6.910 2.310 7.960 2.730 ;
        RECT  6.390 2.130 6.910 2.730 ;
        RECT  5.700 2.310 6.390 2.730 ;
        RECT  5.440 2.290 5.700 2.730 ;
        RECT  4.390 2.310 5.440 2.730 ;
        RECT  4.130 2.115 4.390 2.730 ;
        RECT  3.070 2.310 4.130 2.730 ;
        RECT  2.810 2.190 3.070 2.730 ;
        RECT  1.610 2.310 2.810 2.730 ;
        RECT  0.830 2.220 1.610 2.730 ;
        RECT  0.250 2.310 0.830 2.730 ;
        RECT  0.090 1.550 0.250 2.730 ;
        RECT  0.000 2.310 0.090 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 9.520 2.520 ;
        LAYER M1 ;
        RECT  8.640 0.660 8.760 1.290 ;
        RECT  7.120 0.660 8.640 0.780 ;
        RECT  8.580 1.140 8.640 1.290 ;
        RECT  7.460 1.140 8.580 1.260 ;
        RECT  7.070 0.900 8.470 1.020 ;
        RECT  7.000 0.435 7.120 0.780 ;
        RECT  6.950 0.900 7.070 1.995 ;
        RECT  6.080 0.435 7.000 0.555 ;
        RECT  6.040 1.875 6.950 1.995 ;
        RECT  6.670 0.680 6.790 1.520 ;
        RECT  6.580 1.400 6.670 1.520 ;
        RECT  6.320 1.400 6.580 1.655 ;
        RECT  6.430 0.990 6.550 1.250 ;
        RECT  6.080 1.090 6.430 1.210 ;
        RECT  6.200 1.355 6.320 1.655 ;
        RECT  5.960 0.435 6.080 1.755 ;
        RECT  5.780 1.875 6.040 2.190 ;
        RECT  5.710 0.510 5.960 0.940 ;
        RECT  3.500 1.635 5.960 1.755 ;
        RECT  5.580 1.110 5.820 1.230 ;
        RECT  3.380 1.875 5.780 1.995 ;
        RECT  3.500 0.510 5.710 0.630 ;
        RECT  5.460 0.750 5.580 1.470 ;
        RECT  3.375 0.750 5.460 0.870 ;
        RECT  3.630 1.350 5.460 1.470 ;
        RECT  3.380 1.050 5.140 1.170 ;
        RECT  3.365 1.050 3.380 1.995 ;
        RECT  3.255 0.510 3.375 0.870 ;
        RECT  3.260 1.050 3.365 2.050 ;
        RECT  0.590 1.930 3.260 2.050 ;
        RECT  2.705 0.510 3.255 0.630 ;
        RECT  3.065 1.215 3.140 1.475 ;
        RECT  2.945 0.750 3.065 1.475 ;
        RECT  2.490 0.750 2.945 0.870 ;
        RECT  2.550 1.355 2.945 1.475 ;
        RECT  2.310 1.060 2.825 1.230 ;
        RECT  2.585 0.420 2.705 0.630 ;
        RECT  1.310 0.420 2.585 0.540 ;
        RECT  2.430 1.355 2.550 1.765 ;
        RECT  2.190 0.660 2.310 1.810 ;
        RECT  1.810 0.660 2.190 0.780 ;
        RECT  2.065 1.640 2.190 1.810 ;
        RECT  1.190 0.420 1.310 1.720 ;
        RECT  1.140 1.460 1.190 1.720 ;
        RECT  0.590 1.020 1.070 1.280 ;
        RECT  0.470 0.330 0.590 2.170 ;
    END
END TLATNTSCAX8AD
MACRO TLATNX1AD
    CLASS CORE ;
    FOREIGN TLATNX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 0.655 3.850 1.925 ;
        END
        AntennaDiffArea 0.207 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 1.450 3.105 1.880 ;
        RECT  3.010 0.735 3.065 0.905 ;
        RECT  2.870 0.735 3.010 1.880 ;
        END
        AntennaDiffArea 0.207 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.735 0.210 1.375 ;
        END
        AntennaGateArea 0.068 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.050 1.220 1.310 ;
        RECT  0.910 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.109 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.445 -0.210 3.920 0.210 ;
        RECT  3.275 -0.210 3.445 0.375 ;
        RECT  2.355 -0.210 3.275 0.210 ;
        RECT  2.185 -0.210 2.355 0.795 ;
        RECT  1.075 -0.210 2.185 0.210 ;
        RECT  0.905 -0.210 1.075 0.500 ;
        RECT  0.230 -0.210 0.905 0.210 ;
        RECT  0.110 -0.210 0.230 0.615 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.465 2.310 3.920 2.730 ;
        RECT  3.295 1.450 3.465 2.730 ;
        RECT  2.420 2.310 3.295 2.730 ;
        RECT  2.160 1.750 2.420 2.730 ;
        RECT  1.075 2.310 2.160 2.730 ;
        RECT  0.905 2.030 1.075 2.730 ;
        RECT  0.230 2.310 0.905 2.730 ;
        RECT  0.110 1.850 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  3.440 0.495 3.560 1.270 ;
        RECT  2.690 0.495 3.440 0.615 ;
        RECT  2.690 1.720 2.720 1.980 ;
        RECT  2.570 0.495 2.690 1.980 ;
        RECT  2.070 1.350 2.570 1.610 ;
        RECT  1.950 0.965 2.450 1.225 ;
        RECT  1.830 0.650 1.950 1.870 ;
        RECT  1.680 0.340 1.940 0.500 ;
        RECT  1.680 2.020 1.940 2.180 ;
        RECT  1.510 0.650 1.830 0.770 ;
        RECT  1.510 1.750 1.830 1.870 ;
        RECT  1.315 0.380 1.680 0.500 ;
        RECT  1.390 2.020 1.680 2.140 ;
        RECT  1.470 0.940 1.630 1.060 ;
        RECT  1.390 0.940 1.470 1.600 ;
        RECT  1.350 0.940 1.390 2.140 ;
        RECT  1.270 1.480 1.350 2.140 ;
        RECT  1.195 0.380 1.315 0.740 ;
        RECT  0.615 1.790 1.270 1.910 ;
        RECT  0.710 0.620 1.195 0.740 ;
        RECT  0.710 1.410 0.750 1.670 ;
        RECT  0.590 0.620 0.710 1.670 ;
        RECT  0.470 0.380 0.670 0.500 ;
        RECT  0.470 1.790 0.615 2.065 ;
        RECT  0.445 0.380 0.470 2.065 ;
        RECT  0.350 0.380 0.445 1.910 ;
    END
END TLATNX1AD
MACRO TLATNX2AD
    CLASS CORE ;
    FOREIGN TLATNX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 0.330 3.850 2.190 ;
        END
        AntennaDiffArea 0.368 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 1.455 3.105 2.145 ;
        RECT  3.010 0.735 3.065 0.905 ;
        RECT  2.870 0.735 3.010 2.145 ;
        END
        AntennaDiffArea 0.368 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.735 0.210 1.375 ;
        END
        AntennaGateArea 0.067 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.010 1.220 1.270 ;
        RECT  0.910 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.146 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.445 -0.210 3.920 0.210 ;
        RECT  3.275 -0.210 3.445 0.375 ;
        RECT  2.355 -0.210 3.275 0.210 ;
        RECT  2.185 -0.210 2.355 0.815 ;
        RECT  1.075 -0.210 2.185 0.210 ;
        RECT  0.905 -0.210 1.075 0.475 ;
        RECT  0.230 -0.210 0.905 0.210 ;
        RECT  0.110 -0.210 0.230 0.570 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.465 2.310 3.920 2.730 ;
        RECT  3.295 1.455 3.465 2.730 ;
        RECT  2.420 2.310 3.295 2.730 ;
        RECT  2.160 1.750 2.420 2.730 ;
        RECT  1.075 2.310 2.160 2.730 ;
        RECT  0.905 2.030 1.075 2.730 ;
        RECT  0.230 2.310 0.905 2.730 ;
        RECT  0.110 1.845 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  3.440 0.495 3.560 1.270 ;
        RECT  2.690 0.495 3.440 0.615 ;
        RECT  2.690 1.730 2.720 1.990 ;
        RECT  2.570 0.495 2.690 1.990 ;
        RECT  2.070 1.350 2.570 1.610 ;
        RECT  1.950 0.965 2.450 1.225 ;
        RECT  1.830 0.670 1.950 1.870 ;
        RECT  1.680 0.350 1.940 0.500 ;
        RECT  1.680 2.020 1.940 2.180 ;
        RECT  1.510 0.670 1.830 0.790 ;
        RECT  1.510 1.750 1.830 1.870 ;
        RECT  1.315 0.380 1.680 0.500 ;
        RECT  1.390 2.020 1.680 2.140 ;
        RECT  1.470 0.950 1.630 1.070 ;
        RECT  1.390 0.950 1.470 1.600 ;
        RECT  1.350 0.950 1.390 2.140 ;
        RECT  1.270 1.480 1.350 2.140 ;
        RECT  1.195 0.380 1.315 0.740 ;
        RECT  0.615 1.790 1.270 1.910 ;
        RECT  0.710 0.620 1.195 0.740 ;
        RECT  0.710 1.370 0.750 1.630 ;
        RECT  0.590 0.620 0.710 1.630 ;
        RECT  0.470 0.380 0.670 0.500 ;
        RECT  0.470 1.790 0.615 2.060 ;
        RECT  0.445 0.380 0.470 2.060 ;
        RECT  0.350 0.380 0.445 1.910 ;
    END
END TLATNX2AD
MACRO TLATNX4AD
    CLASS CORE ;
    FOREIGN TLATNX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 0.720 5.530 1.515 ;
        RECT  5.155 0.720 5.390 0.860 ;
        RECT  5.155 1.375 5.390 1.515 ;
        RECT  4.985 0.385 5.155 0.860 ;
        RECT  4.985 1.375 5.155 2.115 ;
        END
        AntennaDiffArea 0.419 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.660 4.410 2.160 ;
        END
        AntennaDiffArea 0.416 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.020 0.230 1.655 ;
        END
        AntennaGateArea 0.117 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.890 1.120 2.105 1.240 ;
        RECT  1.585 1.120 1.890 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.515 -0.210 5.600 0.210 ;
        RECT  5.345 -0.210 5.515 0.600 ;
        RECT  4.820 -0.210 5.345 0.210 ;
        RECT  4.560 -0.210 4.820 0.300 ;
        RECT  4.060 -0.210 4.560 0.210 ;
        RECT  3.800 -0.210 4.060 0.300 ;
        RECT  3.265 -0.210 3.800 0.210 ;
        RECT  3.125 -0.210 3.265 0.870 ;
        RECT  1.985 -0.210 3.125 0.210 ;
        RECT  1.815 -0.210 1.985 0.520 ;
        RECT  0.635 -0.210 1.815 0.210 ;
        RECT  0.465 -0.210 0.635 0.320 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.515 2.310 5.600 2.730 ;
        RECT  5.345 1.635 5.515 2.730 ;
        RECT  4.785 2.310 5.345 2.730 ;
        RECT  4.615 1.425 4.785 2.730 ;
        RECT  4.065 2.310 4.615 2.730 ;
        RECT  3.895 1.675 4.065 2.730 ;
        RECT  3.340 2.310 3.895 2.730 ;
        RECT  3.170 1.995 3.340 2.730 ;
        RECT  1.975 2.310 3.170 2.730 ;
        RECT  1.805 1.975 1.975 2.730 ;
        RECT  0.680 2.310 1.805 2.730 ;
        RECT  0.420 2.240 0.680 2.730 ;
        RECT  0.000 2.310 0.420 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  4.845 1.055 5.270 1.225 ;
        RECT  4.725 0.420 4.845 1.225 ;
        RECT  4.130 0.420 4.725 0.540 ;
        RECT  4.010 0.420 4.130 1.555 ;
        RECT  3.630 0.550 4.010 0.670 ;
        RECT  3.705 1.435 4.010 1.555 ;
        RECT  3.050 1.080 3.815 1.200 ;
        RECT  3.535 1.435 3.705 1.865 ;
        RECT  3.460 0.550 3.630 0.720 ;
        RECT  3.170 1.435 3.535 1.555 ;
        RECT  3.005 1.080 3.050 2.140 ;
        RECT  2.930 0.680 3.005 2.140 ;
        RECT  2.885 0.680 2.930 1.200 ;
        RECT  2.500 2.020 2.930 2.140 ;
        RECT  2.565 0.680 2.885 0.800 ;
        RECT  2.740 1.385 2.810 1.885 ;
        RECT  2.690 0.960 2.740 1.885 ;
        RECT  2.620 0.960 2.690 1.505 ;
        RECT  2.345 0.960 2.620 1.080 ;
        RECT  2.445 0.640 2.565 0.800 ;
        RECT  2.380 1.200 2.500 1.615 ;
        RECT  2.380 1.735 2.500 2.140 ;
        RECT  1.650 0.640 2.445 0.760 ;
        RECT  0.930 1.495 2.380 1.615 ;
        RECT  1.305 1.735 2.380 1.855 ;
        RECT  2.225 0.880 2.345 1.080 ;
        RECT  1.410 0.880 2.225 1.000 ;
        RECT  1.530 0.390 1.650 0.760 ;
        RECT  1.100 0.390 1.530 0.510 ;
        RECT  1.350 0.880 1.410 1.210 ;
        RECT  1.290 0.630 1.350 1.210 ;
        RECT  1.135 1.735 1.305 1.905 ;
        RECT  1.230 0.630 1.290 1.000 ;
        RECT  0.610 0.630 1.230 0.750 ;
        RECT  0.930 2.070 1.090 2.190 ;
        RECT  0.930 0.870 0.990 0.990 ;
        RECT  0.810 0.870 0.930 2.190 ;
        RECT  0.730 0.870 0.810 0.990 ;
        RECT  0.610 1.140 0.680 1.400 ;
        RECT  0.490 0.630 0.610 1.895 ;
        RECT  0.230 0.630 0.490 0.750 ;
        RECT  0.230 1.775 0.490 1.895 ;
        RECT  0.110 0.490 0.230 0.750 ;
        RECT  0.110 1.775 0.230 2.035 ;
    END
END TLATNX4AD
MACRO TLATNXLAD
    CLASS CORE ;
    FOREIGN TLATNXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 0.690 3.850 1.690 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.010 1.475 3.105 1.645 ;
        RECT  3.010 0.735 3.065 0.905 ;
        RECT  2.870 0.735 3.010 1.645 ;
        END
        AntennaDiffArea 0.138 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.735 0.210 1.375 ;
        END
        AntennaGateArea 0.068 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.050 1.220 1.310 ;
        RECT  0.910 0.865 1.050 1.375 ;
        END
        AntennaGateArea 0.086 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.445 -0.210 3.920 0.210 ;
        RECT  3.275 -0.210 3.445 0.375 ;
        RECT  2.355 -0.210 3.275 0.210 ;
        RECT  2.185 -0.210 2.355 0.795 ;
        RECT  1.075 -0.210 2.185 0.210 ;
        RECT  0.905 -0.210 1.075 0.500 ;
        RECT  0.230 -0.210 0.905 0.210 ;
        RECT  0.110 -0.210 0.230 0.615 ;
        RECT  0.000 -0.210 0.110 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.465 2.310 3.920 2.730 ;
        RECT  3.295 1.475 3.465 2.730 ;
        RECT  2.420 2.310 3.295 2.730 ;
        RECT  2.160 1.740 2.420 2.730 ;
        RECT  1.075 2.310 2.160 2.730 ;
        RECT  0.905 2.030 1.075 2.730 ;
        RECT  0.230 2.310 0.905 2.730 ;
        RECT  0.110 1.850 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  3.440 0.495 3.560 1.270 ;
        RECT  2.690 0.495 3.440 0.615 ;
        RECT  2.690 1.710 2.720 1.970 ;
        RECT  2.570 0.495 2.690 1.970 ;
        RECT  2.070 1.350 2.570 1.610 ;
        RECT  1.950 0.965 2.450 1.225 ;
        RECT  1.830 0.650 1.950 1.860 ;
        RECT  1.680 0.340 1.940 0.500 ;
        RECT  1.680 2.020 1.940 2.170 ;
        RECT  1.510 0.650 1.830 0.770 ;
        RECT  1.510 1.740 1.830 1.860 ;
        RECT  1.315 0.380 1.680 0.500 ;
        RECT  1.390 2.020 1.680 2.140 ;
        RECT  1.470 0.940 1.630 1.060 ;
        RECT  1.390 0.940 1.470 1.600 ;
        RECT  1.350 0.940 1.390 2.140 ;
        RECT  1.270 1.480 1.350 2.140 ;
        RECT  1.195 0.380 1.315 0.740 ;
        RECT  0.615 1.790 1.270 1.910 ;
        RECT  0.710 0.620 1.195 0.740 ;
        RECT  0.710 1.410 0.750 1.670 ;
        RECT  0.590 0.620 0.710 1.670 ;
        RECT  0.470 0.380 0.670 0.500 ;
        RECT  0.470 1.790 0.615 2.065 ;
        RECT  0.445 0.380 0.470 2.065 ;
        RECT  0.350 0.380 0.445 1.910 ;
    END
END TLATNXLAD
MACRO TLATSRX1AD
    CLASS CORE ;
    FOREIGN TLATSRX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.855 0.230 1.375 ;
        END
        AntennaGateArea 0.06 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.660 0.850 3.010 1.110 ;
        END
        AntennaGateArea 0.101 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 0.725 5.530 1.905 ;
        RECT  5.345 0.725 5.390 0.895 ;
        RECT  5.360 1.385 5.390 1.905 ;
        END
        AntennaDiffArea 0.205 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.830 0.420 4.970 1.590 ;
        RECT  4.600 0.420 4.830 0.540 ;
        RECT  4.700 1.330 4.830 1.590 ;
        END
        AntennaDiffArea 0.202 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.860 3.350 1.190 ;
        END
        AntennaGateArea 0.068 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.910 1.655 1.330 ;
        END
        AntennaGateArea 0.097 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.225 -0.210 5.600 0.210 ;
        RECT  4.965 -0.210 5.225 0.300 ;
        RECT  4.310 -0.210 4.965 0.210 ;
        RECT  4.050 -0.210 4.310 0.300 ;
        RECT  3.340 -0.210 4.050 0.210 ;
        RECT  3.080 -0.210 3.340 0.300 ;
        RECT  1.440 -0.210 3.080 0.210 ;
        RECT  1.180 -0.210 1.440 0.310 ;
        RECT  0.230 -0.210 1.180 0.210 ;
        RECT  0.070 -0.210 0.230 0.665 ;
        RECT  0.000 -0.210 0.070 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.180 2.310 5.600 2.730 ;
        RECT  4.920 2.220 5.180 2.730 ;
        RECT  4.220 2.310 4.920 2.730 ;
        RECT  3.960 2.220 4.220 2.730 ;
        RECT  3.280 2.310 3.960 2.730 ;
        RECT  3.020 2.270 3.280 2.730 ;
        RECT  1.690 2.310 3.020 2.730 ;
        RECT  1.430 2.220 1.690 2.730 ;
        RECT  0.380 2.310 1.430 2.730 ;
        RECT  0.120 2.220 0.380 2.730 ;
        RECT  0.000 2.310 0.120 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  5.220 1.030 5.270 1.290 ;
        RECT  5.100 1.030 5.220 2.100 ;
        RECT  4.565 1.980 5.100 2.100 ;
        RECT  4.430 0.735 4.565 2.100 ;
        RECT  4.395 0.735 4.430 0.905 ;
        RECT  3.020 1.980 4.430 2.100 ;
        RECT  4.190 1.040 4.310 1.840 ;
        RECT  0.870 1.720 4.190 1.840 ;
        RECT  3.840 0.370 3.950 1.460 ;
        RECT  3.830 0.370 3.840 1.600 ;
        RECT  3.670 0.370 3.830 0.540 ;
        RECT  3.720 1.340 3.830 1.600 ;
        RECT  3.600 0.960 3.710 1.220 ;
        RECT  2.580 0.420 3.670 0.540 ;
        RECT  3.480 0.670 3.600 1.600 ;
        RECT  2.400 1.480 3.480 1.600 ;
        RECT  2.760 1.980 3.020 2.150 ;
        RECT  2.460 0.420 2.580 0.740 ;
        RECT  2.400 0.890 2.540 1.010 ;
        RECT  2.160 0.620 2.460 0.740 ;
        RECT  2.280 0.890 2.400 1.600 ;
        RECT  1.920 0.380 2.340 0.500 ;
        RECT  1.110 1.480 2.280 1.600 ;
        RECT  1.940 1.980 2.200 2.190 ;
        RECT  2.040 0.620 2.160 1.270 ;
        RECT  1.980 1.010 2.040 1.270 ;
        RECT  0.530 1.980 1.940 2.100 ;
        RECT  1.800 0.380 1.920 0.600 ;
        RECT  1.255 0.480 1.800 0.600 ;
        RECT  1.135 0.480 1.255 0.810 ;
        RECT  0.710 0.690 1.135 0.810 ;
        RECT  0.990 1.095 1.110 1.600 ;
        RECT  0.950 1.095 0.990 1.215 ;
        RECT  0.710 0.380 0.970 0.570 ;
        RECT  0.830 0.955 0.950 1.215 ;
        RECT  0.750 1.335 0.870 1.840 ;
        RECT  0.710 1.335 0.750 1.455 ;
        RECT  0.470 0.450 0.710 0.570 ;
        RECT  0.590 0.690 0.710 1.455 ;
        RECT  0.470 1.600 0.530 2.100 ;
        RECT  0.350 0.450 0.470 2.100 ;
    END
END TLATSRX1AD
MACRO TLATSRX2AD
    CLASS CORE ;
    FOREIGN TLATSRX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.085 0.230 1.655 ;
        END
        AntennaGateArea 0.091 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.810 0.865 3.010 1.235 ;
        END
        AntennaGateArea 0.152 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.930 0.365 6.090 2.190 ;
        END
        AntennaDiffArea 0.373 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.250 0.410 5.305 0.840 ;
        RECT  5.210 0.410 5.250 1.095 ;
        RECT  5.050 0.410 5.210 1.850 ;
        END
        AntennaDiffArea 0.373 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.070 3.560 1.330 ;
        RECT  3.150 0.865 3.290 1.330 ;
        END
        AntennaGateArea 0.067 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.425 0.910 1.690 1.330 ;
        END
        AntennaGateArea 0.139 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.695 -0.210 6.160 0.210 ;
        RECT  5.525 -0.210 5.695 0.830 ;
        RECT  4.620 -0.210 5.525 0.210 ;
        RECT  4.360 -0.210 4.620 0.660 ;
        RECT  3.500 -0.210 4.360 0.210 ;
        RECT  3.240 -0.210 3.500 0.300 ;
        RECT  1.520 -0.210 3.240 0.210 ;
        RECT  1.260 -0.210 1.520 0.300 ;
        RECT  0.230 -0.210 1.260 0.210 ;
        RECT  0.070 -0.210 0.230 0.810 ;
        RECT  0.000 -0.210 0.070 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.730 2.310 6.160 2.730 ;
        RECT  5.570 1.800 5.730 2.730 ;
        RECT  4.620 2.310 5.570 2.730 ;
        RECT  4.360 2.220 4.620 2.730 ;
        RECT  3.580 2.310 4.360 2.730 ;
        RECT  3.320 2.220 3.580 2.730 ;
        RECT  1.840 2.310 3.320 2.730 ;
        RECT  1.580 2.170 1.840 2.730 ;
        RECT  0.230 2.310 1.580 2.730 ;
        RECT  0.070 1.820 0.230 2.730 ;
        RECT  0.000 2.310 0.070 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.640 0.995 5.760 1.465 ;
        RECT  5.450 1.345 5.640 1.465 ;
        RECT  5.330 1.345 5.450 2.100 ;
        RECT  4.860 1.980 5.330 2.100 ;
        RECT  4.860 0.585 4.930 0.845 ;
        RECT  4.740 0.585 4.860 2.100 ;
        RECT  3.200 1.980 4.740 2.100 ;
        RECT  4.500 1.040 4.620 1.860 ;
        RECT  3.440 1.740 4.500 1.860 ;
        RECT  4.260 0.785 4.380 1.480 ;
        RECT  4.170 0.785 4.260 0.905 ;
        RECT  4.170 1.360 4.260 1.480 ;
        RECT  4.050 0.420 4.170 0.905 ;
        RECT  4.050 1.360 4.170 1.620 ;
        RECT  3.900 1.025 4.140 1.195 ;
        RECT  2.720 0.420 4.050 0.540 ;
        RECT  3.780 0.705 3.900 1.620 ;
        RECT  3.665 0.705 3.780 0.875 ;
        RECT  3.640 1.450 3.780 1.620 ;
        RECT  2.615 1.450 3.640 1.570 ;
        RECT  3.320 1.690 3.440 1.860 ;
        RECT  0.950 1.690 3.320 1.810 ;
        RECT  3.080 1.930 3.200 2.190 ;
        RECT  2.780 1.930 2.900 2.190 ;
        RECT  0.660 1.930 2.780 2.050 ;
        RECT  2.600 0.420 2.720 0.765 ;
        RECT  2.615 0.900 2.685 1.020 ;
        RECT  2.495 0.900 2.615 1.570 ;
        RECT  2.240 0.645 2.600 0.765 ;
        RECT  2.425 0.900 2.495 1.020 ;
        RECT  1.190 1.450 2.495 1.570 ;
        RECT  1.775 0.405 2.480 0.525 ;
        RECT  2.240 1.155 2.375 1.300 ;
        RECT  2.115 0.645 2.240 1.300 ;
        RECT  1.655 0.405 1.775 0.720 ;
        RECT  0.990 0.600 1.655 0.720 ;
        RECT  1.070 1.135 1.190 1.570 ;
        RECT  0.840 1.135 1.070 1.255 ;
        RECT  0.870 0.600 0.990 0.980 ;
        RECT  0.830 1.510 0.950 1.810 ;
        RECT  0.710 0.860 0.870 0.980 ;
        RECT  0.660 0.330 0.865 0.450 ;
        RECT  0.710 1.510 0.830 1.690 ;
        RECT  0.590 0.860 0.710 1.690 ;
        RECT  0.540 0.330 0.660 0.740 ;
        RECT  0.470 1.850 0.660 2.050 ;
        RECT  0.470 0.620 0.540 0.740 ;
        RECT  0.350 0.620 0.470 2.050 ;
    END
END TLATSRX2AD
MACRO TLATSRX4AD
    CLASS CORE ;
    FOREIGN TLATSRX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.000 0.390 1.260 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.790 0.825 4.910 1.300 ;
        RECT  4.175 1.180 4.790 1.300 ;
        RECT  3.765 1.180 4.175 1.330 ;
        RECT  3.645 0.910 3.765 1.330 ;
        RECT  2.530 0.910 3.645 1.030 ;
        RECT  2.270 0.910 2.530 1.070 ;
        END
        AntennaGateArea 0.259 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.330 0.405 8.485 0.865 ;
        RECT  8.330 1.330 8.470 1.590 ;
        RECT  8.315 0.405 8.330 1.590 ;
        RECT  8.190 0.725 8.315 1.590 ;
        END
        AntennaDiffArea 0.462 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.630 0.410 7.770 1.590 ;
        RECT  7.555 0.410 7.630 0.840 ;
        RECT  7.555 1.420 7.630 1.590 ;
        END
        AntennaDiffArea 0.454 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  5.390 0.865 5.550 1.290 ;
        END
        AntennaGateArea 0.1 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.620 1.180 2.880 1.375 ;
        RECT  2.110 1.255 2.620 1.375 ;
        RECT  1.890 1.200 2.110 1.375 ;
        RECT  1.470 1.145 1.890 1.375 ;
        END
        AntennaGateArea 0.291 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.855 -0.210 8.960 0.210 ;
        RECT  8.695 -0.210 8.855 0.860 ;
        RECT  8.105 -0.210 8.695 0.210 ;
        RECT  7.935 -0.210 8.105 0.605 ;
        RECT  7.355 -0.210 7.935 0.210 ;
        RECT  7.355 0.435 7.400 0.815 ;
        RECT  7.185 -0.210 7.355 0.840 ;
        RECT  6.660 -0.210 7.185 0.210 ;
        RECT  7.140 0.435 7.185 0.815 ;
        RECT  6.400 -0.210 6.660 0.585 ;
        RECT  5.500 -0.210 6.400 0.210 ;
        RECT  5.240 -0.210 5.500 0.415 ;
        RECT  3.425 -0.210 5.240 0.210 ;
        RECT  2.905 -0.210 3.425 0.300 ;
        RECT  1.430 -0.210 2.905 0.210 ;
        RECT  1.170 -0.210 1.430 0.500 ;
        RECT  0.680 -0.210 1.170 0.210 ;
        RECT  0.420 -0.210 0.680 0.505 ;
        RECT  0.000 -0.210 0.420 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  8.855 2.310 8.960 2.730 ;
        RECT  8.675 1.950 8.855 2.730 ;
        RECT  8.120 2.310 8.675 2.730 ;
        RECT  7.920 1.950 8.120 2.730 ;
        RECT  7.370 2.310 7.920 2.730 ;
        RECT  7.170 1.950 7.370 2.730 ;
        RECT  6.660 2.310 7.170 2.730 ;
        RECT  6.400 2.220 6.660 2.730 ;
        RECT  5.660 2.310 6.400 2.730 ;
        RECT  5.400 2.255 5.660 2.730 ;
        RECT  3.990 2.310 5.400 2.730 ;
        RECT  3.730 2.220 3.990 2.730 ;
        RECT  1.990 2.310 3.730 2.730 ;
        RECT  1.730 2.220 1.990 2.730 ;
        RECT  0.625 2.310 1.730 2.730 ;
        RECT  0.455 2.105 0.625 2.730 ;
        RECT  0.000 2.310 0.455 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 8.960 2.520 ;
        LAYER M1 ;
        RECT  8.590 1.030 8.710 1.830 ;
        RECT  8.450 1.030 8.590 1.190 ;
        RECT  6.970 1.710 8.590 1.830 ;
        RECT  6.850 0.535 6.970 2.100 ;
        RECT  5.280 1.980 6.850 2.100 ;
        RECT  6.590 1.005 6.710 1.860 ;
        RECT  5.530 1.740 6.590 1.860 ;
        RECT  6.350 0.705 6.470 1.480 ;
        RECT  6.210 0.705 6.350 0.830 ;
        RECT  6.210 1.360 6.350 1.480 ;
        RECT  5.940 0.980 6.230 1.240 ;
        RECT  6.090 0.535 6.210 0.830 ;
        RECT  6.090 1.360 6.210 1.620 ;
        RECT  4.660 0.535 6.090 0.655 ;
        RECT  5.815 0.785 5.940 1.595 ;
        RECT  5.670 0.785 5.815 0.905 ;
        RECT  5.670 1.450 5.815 1.595 ;
        RECT  4.750 1.450 5.670 1.570 ;
        RECT  5.410 1.690 5.530 1.860 ;
        RECT  4.970 1.690 5.410 1.810 ;
        RECT  5.160 1.930 5.280 2.190 ;
        RECT  4.750 1.980 5.010 2.190 ;
        RECT  4.850 1.690 4.970 1.860 ;
        RECT  1.110 1.740 4.850 1.860 ;
        RECT  4.630 1.450 4.750 1.620 ;
        RECT  3.550 1.980 4.750 2.100 ;
        RECT  4.540 0.535 4.660 1.060 ;
        RECT  3.280 1.500 4.630 1.620 ;
        RECT  4.120 0.920 4.540 1.060 ;
        RECT  4.240 0.430 4.360 0.690 ;
        RECT  1.850 0.430 4.240 0.550 ;
        RECT  3.995 0.670 4.120 1.060 ;
        RECT  2.125 0.670 3.995 0.790 ;
        RECT  3.290 1.980 3.550 2.190 ;
        RECT  2.810 1.980 3.290 2.100 ;
        RECT  3.020 1.190 3.280 1.620 ;
        RECT  1.350 1.500 3.020 1.620 ;
        RECT  2.550 1.980 2.810 2.190 ;
        RECT  0.865 1.980 2.550 2.100 ;
        RECT  1.990 0.670 2.125 0.990 ;
        RECT  1.580 0.860 1.990 0.990 ;
        RECT  1.700 0.430 1.850 0.740 ;
        RECT  1.000 0.620 1.700 0.740 ;
        RECT  1.230 1.225 1.350 1.620 ;
        RECT  1.190 1.225 1.230 1.355 ;
        RECT  1.070 1.095 1.190 1.355 ;
        RECT  0.990 1.480 1.110 1.860 ;
        RECT  0.950 0.395 1.000 0.740 ;
        RECT  0.950 1.480 0.990 1.740 ;
        RECT  0.830 0.395 0.950 1.740 ;
        RECT  0.745 1.860 0.865 2.100 ;
        RECT  0.630 1.860 0.745 1.985 ;
        RECT  0.630 0.980 0.710 1.240 ;
        RECT  0.510 0.625 0.630 1.985 ;
        RECT  0.240 0.625 0.510 0.745 ;
        RECT  0.265 1.860 0.510 1.985 ;
        RECT  0.095 1.555 0.265 1.985 ;
        RECT  0.080 0.485 0.240 0.745 ;
    END
END TLATSRX4AD
MACRO TLATSRXLAD
    CLASS CORE ;
    FOREIGN TLATSRXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.855 0.230 1.375 ;
        RECT  0.070 1.145 0.090 1.375 ;
        END
        AntennaGateArea 0.051 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.680 0.850 3.010 1.110 ;
        END
        AntennaGateArea 0.085 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 0.590 5.530 1.635 ;
        RECT  5.330 0.590 5.390 0.850 ;
        RECT  5.345 1.465 5.390 1.635 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 0.865 4.970 1.375 ;
        RECT  4.770 0.420 4.890 1.545 ;
        RECT  4.610 0.420 4.770 0.540 ;
        RECT  4.675 1.375 4.770 1.545 ;
        END
        AntennaDiffArea 0.157 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  3.150 0.860 3.350 1.240 ;
        END
        AntennaGateArea 0.068 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.415 0.910 1.655 1.330 ;
        END
        AntennaGateArea 0.075 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.215 -0.210 5.600 0.210 ;
        RECT  4.955 -0.210 5.215 0.300 ;
        RECT  4.310 -0.210 4.955 0.210 ;
        RECT  4.050 -0.210 4.310 0.300 ;
        RECT  3.340 -0.210 4.050 0.210 ;
        RECT  3.080 -0.210 3.340 0.300 ;
        RECT  1.440 -0.210 3.080 0.210 ;
        RECT  1.180 -0.210 1.440 0.300 ;
        RECT  0.230 -0.210 1.180 0.210 ;
        RECT  0.070 -0.210 0.230 0.640 ;
        RECT  0.000 -0.210 0.070 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.180 2.310 5.600 2.730 ;
        RECT  4.920 2.220 5.180 2.730 ;
        RECT  4.220 2.310 4.920 2.730 ;
        RECT  3.960 2.220 4.220 2.730 ;
        RECT  3.390 2.310 3.960 2.730 ;
        RECT  3.130 2.220 3.390 2.730 ;
        RECT  1.690 2.310 3.130 2.730 ;
        RECT  1.430 2.220 1.690 2.730 ;
        RECT  0.380 2.310 1.430 2.730 ;
        RECT  0.120 2.220 0.380 2.730 ;
        RECT  0.000 2.310 0.120 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  5.220 1.010 5.270 1.270 ;
        RECT  5.100 1.010 5.220 2.100 ;
        RECT  4.555 1.980 5.100 2.100 ;
        RECT  4.555 0.735 4.565 0.905 ;
        RECT  4.430 0.735 4.555 2.100 ;
        RECT  4.395 0.735 4.430 0.905 ;
        RECT  3.020 1.980 4.430 2.100 ;
        RECT  4.190 1.050 4.310 1.840 ;
        RECT  0.870 1.720 4.190 1.840 ;
        RECT  3.830 0.370 3.950 1.600 ;
        RECT  3.670 0.370 3.830 0.540 ;
        RECT  3.720 1.340 3.830 1.600 ;
        RECT  3.600 0.960 3.710 1.220 ;
        RECT  2.580 0.420 3.670 0.540 ;
        RECT  3.480 0.670 3.600 1.600 ;
        RECT  2.400 1.480 3.480 1.600 ;
        RECT  2.760 1.980 3.020 2.150 ;
        RECT  2.460 0.420 2.580 0.740 ;
        RECT  2.400 0.890 2.540 1.010 ;
        RECT  2.160 0.620 2.460 0.740 ;
        RECT  2.280 0.890 2.400 1.600 ;
        RECT  1.920 0.380 2.340 0.500 ;
        RECT  1.110 1.480 2.280 1.600 ;
        RECT  1.940 1.980 2.200 2.190 ;
        RECT  2.040 0.620 2.160 1.270 ;
        RECT  1.980 1.010 2.040 1.270 ;
        RECT  0.530 1.980 1.940 2.100 ;
        RECT  1.800 0.380 1.920 0.600 ;
        RECT  1.190 0.480 1.800 0.600 ;
        RECT  1.070 0.480 1.190 0.810 ;
        RECT  0.990 1.095 1.110 1.600 ;
        RECT  0.710 0.690 1.070 0.810 ;
        RECT  0.950 1.095 0.990 1.215 ;
        RECT  0.690 0.330 0.950 0.570 ;
        RECT  0.830 0.955 0.950 1.215 ;
        RECT  0.750 1.335 0.870 1.840 ;
        RECT  0.710 1.335 0.750 1.455 ;
        RECT  0.590 0.690 0.710 1.455 ;
        RECT  0.470 0.450 0.690 0.570 ;
        RECT  0.470 1.600 0.530 2.100 ;
        RECT  0.350 0.450 0.470 2.100 ;
    END
END TLATSRXLAD
MACRO TLATX1AD
    CLASS CORE ;
    FOREIGN TLATX1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 0.690 3.570 1.925 ;
        RECT  3.385 0.690 3.430 0.860 ;
        RECT  3.400 1.405 3.430 1.925 ;
        END
        AntennaDiffArea 0.207 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.425 3.010 1.655 ;
        RECT  2.740 0.690 2.860 1.655 ;
        END
        AntennaDiffArea 0.178 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.210 1.370 ;
        END
        AntennaGateArea 0.049 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.230 1.170 1.655 ;
        END
        AntennaGateArea 0.109 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.265 -0.210 3.640 0.210 ;
        RECT  3.095 -0.210 3.265 0.330 ;
        RECT  2.255 -0.210 3.095 0.210 ;
        RECT  2.085 -0.210 2.255 0.330 ;
        RECT  0.960 -0.210 2.085 0.210 ;
        RECT  0.530 -0.210 0.960 0.310 ;
        RECT  0.000 -0.210 0.530 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.175 2.310 3.640 2.730 ;
        RECT  3.005 2.195 3.175 2.730 ;
        RECT  2.305 2.310 3.005 2.730 ;
        RECT  2.135 2.260 2.305 2.730 ;
        RECT  1.080 2.310 2.135 2.730 ;
        RECT  0.820 2.020 1.080 2.730 ;
        RECT  0.265 2.310 0.820 2.730 ;
        RECT  0.095 1.525 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  3.190 1.010 3.310 1.270 ;
        RECT  3.100 1.010 3.190 1.130 ;
        RECT  2.980 0.450 3.100 1.130 ;
        RECT  2.635 0.450 2.980 0.570 ;
        RECT  2.465 0.355 2.635 0.570 ;
        RECT  2.500 1.090 2.620 1.935 ;
        RECT  2.310 1.090 2.500 1.210 ;
        RECT  2.445 1.765 2.500 1.935 ;
        RECT  2.310 0.450 2.465 0.570 ;
        RECT  2.260 1.330 2.380 1.590 ;
        RECT  2.190 0.450 2.310 1.210 ;
        RECT  2.070 1.470 2.260 1.590 ;
        RECT  1.950 0.510 2.070 2.140 ;
        RECT  1.430 0.510 1.950 0.630 ;
        RECT  1.435 2.020 1.950 2.140 ;
        RECT  1.710 0.750 1.830 1.240 ;
        RECT  1.690 1.640 1.810 1.900 ;
        RECT  1.295 0.750 1.710 0.870 ;
        RECT  1.430 1.780 1.690 1.900 ;
        RECT  1.430 0.990 1.570 1.140 ;
        RECT  1.310 0.990 1.430 1.900 ;
        RECT  1.055 0.990 1.310 1.110 ;
        RECT  0.675 1.780 1.310 1.900 ;
        RECT  1.175 0.430 1.295 0.870 ;
        RECT  0.450 0.430 1.175 0.550 ;
        RECT  0.935 0.810 1.055 1.110 ;
        RECT  0.695 0.810 0.935 0.930 ;
        RECT  0.670 1.125 0.790 1.660 ;
        RECT  0.575 0.670 0.695 0.930 ;
        RECT  0.505 1.780 0.675 2.125 ;
        RECT  0.450 1.125 0.670 1.245 ;
        RECT  0.410 1.540 0.670 1.660 ;
        RECT  0.330 0.430 0.450 1.245 ;
        RECT  0.265 0.430 0.330 0.550 ;
        RECT  0.095 0.375 0.265 0.550 ;
    END
END TLATX1AD
MACRO TLATX2AD
    CLASS CORE ;
    FOREIGN TLATX2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.680 0.330 3.850 2.190 ;
        END
        AntennaDiffArea 0.368 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.080 0.865 3.290 1.095 ;
        RECT  2.920 0.680 3.080 2.190 ;
        END
        AntennaDiffArea 0.368 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.735 0.210 1.375 ;
        END
        AntennaGateArea 0.064 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.100 0.865 1.220 1.290 ;
        RECT  0.910 0.865 1.100 1.095 ;
        END
        AntennaGateArea 0.15 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.490 -0.210 3.920 0.210 ;
        RECT  3.230 -0.210 3.490 0.320 ;
        RECT  2.440 -0.210 3.230 0.210 ;
        RECT  2.180 -0.210 2.440 0.330 ;
        RECT  1.070 -0.210 2.180 0.210 ;
        RECT  0.810 -0.210 1.070 0.310 ;
        RECT  0.230 -0.210 0.810 0.210 ;
        RECT  0.070 -0.210 0.230 0.555 ;
        RECT  0.000 -0.210 0.070 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.465 2.310 3.920 2.730 ;
        RECT  3.295 1.455 3.465 2.730 ;
        RECT  2.395 2.310 3.295 2.730 ;
        RECT  2.215 1.755 2.395 2.730 ;
        RECT  1.095 2.310 2.215 2.730 ;
        RECT  0.925 1.995 1.095 2.730 ;
        RECT  0.230 2.310 0.925 2.730 ;
        RECT  0.110 1.910 0.230 2.730 ;
        RECT  0.000 2.310 0.110 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.920 2.520 ;
        LAYER M1 ;
        RECT  3.440 0.440 3.560 1.270 ;
        RECT  2.800 0.440 3.440 0.560 ;
        RECT  2.730 0.440 2.800 1.430 ;
        RECT  2.680 0.440 2.730 1.985 ;
        RECT  2.570 0.610 2.680 0.870 ;
        RECT  2.610 1.310 2.680 1.985 ;
        RECT  2.200 1.310 2.610 1.430 ;
        RECT  1.870 1.040 2.560 1.160 ;
        RECT  2.080 1.310 2.200 1.570 ;
        RECT  1.690 2.020 1.950 2.190 ;
        RECT  1.680 0.330 1.940 0.500 ;
        RECT  1.750 0.690 1.870 1.885 ;
        RECT  1.510 0.690 1.750 0.810 ;
        RECT  1.555 1.715 1.750 1.885 ;
        RECT  1.380 2.020 1.690 2.140 ;
        RECT  1.380 0.380 1.680 0.500 ;
        RECT  1.460 1.000 1.630 1.120 ;
        RECT  1.380 1.000 1.460 1.610 ;
        RECT  1.260 0.380 1.380 0.550 ;
        RECT  1.340 1.000 1.380 2.140 ;
        RECT  1.260 1.490 1.340 2.140 ;
        RECT  0.615 0.430 1.260 0.550 ;
        RECT  0.760 1.490 1.260 1.610 ;
        RECT  0.640 0.670 0.760 1.725 ;
        RECT  0.470 0.340 0.615 0.550 ;
        RECT  0.470 1.960 0.615 2.130 ;
        RECT  0.350 0.340 0.470 2.130 ;
    END
END TLATX2AD
MACRO TLATX4AD
    CLASS CORE ;
    FOREIGN TLATX4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 0.720 5.530 1.515 ;
        RECT  5.155 0.720 5.390 0.860 ;
        RECT  5.145 1.375 5.390 1.515 ;
        RECT  4.985 0.360 5.155 0.860 ;
        RECT  4.975 1.375 5.145 2.170 ;
        END
        AntennaDiffArea 0.429 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 0.690 4.425 2.170 ;
        END
        AntennaDiffArea 0.416 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.055 0.370 1.225 ;
        RECT  0.070 1.055 0.210 1.375 ;
        END
        AntennaGateArea 0.108 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.100 2.070 1.375 ;
        END
        AntennaGateArea 0.314 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.515 -0.210 5.600 0.210 ;
        RECT  5.345 -0.210 5.515 0.600 ;
        RECT  4.775 -0.210 5.345 0.210 ;
        RECT  4.605 -0.210 4.775 0.330 ;
        RECT  4.015 -0.210 4.605 0.210 ;
        RECT  3.845 -0.210 4.015 0.330 ;
        RECT  3.290 -0.210 3.845 0.210 ;
        RECT  3.170 -0.210 3.290 0.775 ;
        RECT  1.985 -0.210 3.170 0.210 ;
        RECT  1.815 -0.210 1.985 0.500 ;
        RECT  0.615 -0.210 1.815 0.210 ;
        RECT  0.445 -0.210 0.615 0.675 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  5.515 2.310 5.600 2.730 ;
        RECT  5.345 1.635 5.515 2.730 ;
        RECT  4.785 2.310 5.345 2.730 ;
        RECT  4.615 1.480 4.785 2.730 ;
        RECT  4.065 2.310 4.615 2.730 ;
        RECT  3.895 1.675 4.065 2.730 ;
        RECT  3.290 2.310 3.895 2.730 ;
        RECT  3.170 1.865 3.290 2.730 ;
        RECT  1.975 2.310 3.170 2.730 ;
        RECT  1.805 1.975 1.975 2.730 ;
        RECT  0.635 2.310 1.805 2.730 ;
        RECT  0.465 1.905 0.635 2.730 ;
        RECT  0.000 2.310 0.465 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.600 2.520 ;
        LAYER M1 ;
        RECT  4.800 1.080 5.270 1.200 ;
        RECT  4.680 0.450 4.800 1.200 ;
        RECT  4.130 0.450 4.680 0.570 ;
        RECT  4.010 0.450 4.130 1.550 ;
        RECT  3.505 0.560 4.010 0.730 ;
        RECT  3.685 1.430 4.010 1.550 ;
        RECT  3.050 1.075 3.890 1.195 ;
        RECT  3.515 1.430 3.685 1.860 ;
        RECT  3.340 1.430 3.515 1.550 ;
        RECT  3.170 1.380 3.340 1.550 ;
        RECT  2.930 0.620 3.050 2.055 ;
        RECT  2.705 0.620 2.930 0.740 ;
        RECT  2.500 1.935 2.930 2.055 ;
        RECT  2.690 0.970 2.810 1.815 ;
        RECT  2.445 0.330 2.705 0.740 ;
        RECT  2.375 0.970 2.690 1.090 ;
        RECT  2.430 1.270 2.570 1.390 ;
        RECT  2.380 1.735 2.500 2.055 ;
        RECT  1.360 0.620 2.445 0.740 ;
        RECT  2.310 1.270 2.430 1.615 ;
        RECT  1.535 1.735 2.380 1.855 ;
        RECT  2.255 0.860 2.375 1.090 ;
        RECT  1.255 1.495 2.310 1.615 ;
        RECT  1.480 0.860 2.255 0.980 ;
        RECT  1.415 1.735 1.535 2.025 ;
        RECT  1.360 0.860 1.480 1.090 ;
        RECT  1.280 1.905 1.415 2.025 ;
        RECT  1.240 0.330 1.360 0.740 ;
        RECT  0.970 0.970 1.360 1.090 ;
        RECT  1.160 1.905 1.280 2.165 ;
        RECT  1.135 1.495 1.255 1.785 ;
        RECT  1.100 0.330 1.240 0.450 ;
        RECT  1.015 1.665 1.135 1.785 ;
        RECT  0.970 1.375 1.015 1.545 ;
        RECT  0.755 1.665 1.015 2.190 ;
        RECT  0.830 0.570 0.970 1.545 ;
        RECT  0.610 1.665 0.755 1.785 ;
        RECT  0.610 1.000 0.680 1.260 ;
        RECT  0.490 0.815 0.610 1.785 ;
        RECT  0.255 0.815 0.490 0.935 ;
        RECT  0.255 1.665 0.490 1.785 ;
        RECT  0.085 0.520 0.255 0.935 ;
        RECT  0.085 1.495 0.255 1.925 ;
    END
END TLATX4AD
MACRO TLATXLAD
    CLASS CORE ;
    FOREIGN TLATXLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.640 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.430 0.735 3.570 1.645 ;
        RECT  3.385 0.735 3.430 0.905 ;
        RECT  3.385 1.475 3.430 1.645 ;
        END
        AntennaDiffArea 0.138 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.425 3.010 1.655 ;
        RECT  2.740 0.690 2.860 1.655 ;
        END
        AntennaDiffArea 0.134 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.865 0.210 1.370 ;
        END
        AntennaGateArea 0.048 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.230 1.170 1.655 ;
        END
        AntennaGateArea 0.086 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.265 -0.210 3.640 0.210 ;
        RECT  3.095 -0.210 3.265 0.330 ;
        RECT  2.255 -0.210 3.095 0.210 ;
        RECT  2.085 -0.210 2.255 0.330 ;
        RECT  0.960 -0.210 2.085 0.210 ;
        RECT  0.530 -0.210 0.960 0.310 ;
        RECT  0.000 -0.210 0.530 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  3.175 2.310 3.640 2.730 ;
        RECT  3.005 2.005 3.175 2.730 ;
        RECT  2.305 2.310 3.005 2.730 ;
        RECT  2.135 2.260 2.305 2.730 ;
        RECT  1.080 2.310 2.135 2.730 ;
        RECT  0.820 2.020 1.080 2.730 ;
        RECT  0.265 2.310 0.820 2.730 ;
        RECT  0.095 1.515 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.640 2.520 ;
        LAYER M1 ;
        RECT  3.190 1.010 3.310 1.270 ;
        RECT  3.100 1.010 3.190 1.130 ;
        RECT  2.980 0.450 3.100 1.130 ;
        RECT  2.635 0.450 2.980 0.570 ;
        RECT  2.465 0.355 2.635 0.570 ;
        RECT  2.500 1.090 2.620 1.935 ;
        RECT  2.310 1.090 2.500 1.210 ;
        RECT  2.445 1.765 2.500 1.935 ;
        RECT  2.310 0.450 2.465 0.570 ;
        RECT  2.260 1.330 2.380 1.590 ;
        RECT  2.190 0.450 2.310 1.210 ;
        RECT  2.070 1.470 2.260 1.590 ;
        RECT  1.950 0.510 2.070 2.140 ;
        RECT  1.430 0.510 1.950 0.630 ;
        RECT  1.435 2.020 1.950 2.140 ;
        RECT  1.710 0.750 1.830 1.240 ;
        RECT  1.690 1.640 1.810 1.900 ;
        RECT  1.295 0.750 1.710 0.870 ;
        RECT  1.430 1.780 1.690 1.900 ;
        RECT  1.430 0.990 1.570 1.110 ;
        RECT  1.310 0.990 1.430 1.900 ;
        RECT  1.055 0.990 1.310 1.110 ;
        RECT  0.675 1.780 1.310 1.900 ;
        RECT  1.175 0.430 1.295 0.870 ;
        RECT  0.450 0.430 1.175 0.550 ;
        RECT  0.935 0.810 1.055 1.110 ;
        RECT  0.695 0.810 0.935 0.930 ;
        RECT  0.670 1.125 0.790 1.660 ;
        RECT  0.575 0.670 0.695 0.930 ;
        RECT  0.505 1.780 0.675 2.125 ;
        RECT  0.450 1.125 0.670 1.245 ;
        RECT  0.410 1.540 0.670 1.660 ;
        RECT  0.330 0.430 0.450 1.245 ;
        RECT  0.265 0.430 0.330 0.550 ;
        RECT  0.095 0.375 0.265 0.550 ;
    END
END TLATXLAD
MACRO XNOR2X1AD
    CLASS CORE ;
    FOREIGN XNOR2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.350 1.655 0.490 ;
        RECT  1.430 0.350 1.550 1.850 ;
        RECT  1.145 0.350 1.430 0.680 ;
        RECT  1.200 1.730 1.430 1.850 ;
        END
        AntennaDiffArea 0.16 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 0.865 0.770 1.105 ;
        END
        AntennaGateArea 0.088 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.200 1.705 0.490 2.170 ;
        END
        AntennaGateArea 0.1074 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.090 -0.210 2.240 0.210 ;
        RECT  1.970 -0.210 2.090 0.400 ;
        RECT  0.645 -0.210 1.970 0.210 ;
        RECT  0.475 -0.210 0.645 0.705 ;
        RECT  0.000 -0.210 0.475 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 2.310 2.240 2.730 ;
        RECT  1.880 2.220 2.140 2.730 ;
        RECT  0.730 2.310 1.880 2.730 ;
        RECT  0.610 1.465 0.730 2.730 ;
        RECT  0.420 1.465 0.610 1.585 ;
        RECT  0.000 2.310 0.610 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.920 1.020 2.040 2.090 ;
        RECT  1.010 1.970 1.920 2.090 ;
        RECT  1.670 0.670 1.790 1.850 ;
        RECT  1.190 0.800 1.310 1.610 ;
        RECT  1.025 0.800 1.190 0.920 ;
        RECT  1.010 1.490 1.190 1.610 ;
        RECT  0.950 1.040 1.070 1.345 ;
        RECT  0.890 0.560 1.025 0.920 ;
        RECT  0.890 1.490 1.010 2.090 ;
        RECT  0.265 1.225 0.950 1.345 ;
        RECT  0.855 0.560 0.890 0.730 ;
        RECT  0.225 0.625 0.265 0.795 ;
        RECT  0.225 1.225 0.265 1.555 ;
        RECT  0.095 0.625 0.225 1.555 ;
    END
END XNOR2X1AD
MACRO XNOR2X2AD
    CLASS CORE ;
    FOREIGN XNOR2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.080 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.345 2.495 1.895 ;
        RECT  2.280 0.345 2.310 0.775 ;
        END
        AntennaDiffArea 0.387 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.240 1.020 0.345 1.280 ;
        RECT  0.070 0.865 0.240 1.375 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 0.845 1.610 1.380 ;
        END
        AntennaGateArea 0.1927 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.365 -0.210 3.080 0.210 ;
        RECT  1.180 -0.210 1.365 0.675 ;
        RECT  0.265 -0.210 1.180 0.210 ;
        RECT  0.095 -0.210 0.265 0.675 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  1.465 2.310 3.080 2.730 ;
        RECT  1.205 2.220 1.465 2.730 ;
        RECT  0.270 2.310 1.205 2.730 ;
        RECT  0.100 1.585 0.270 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 3.080 2.520 ;
        LAYER M1 ;
        RECT  2.705 0.345 2.875 2.140 ;
        RECT  2.650 0.345 2.705 0.775 ;
        RECT  1.885 2.015 2.705 2.140 ;
        RECT  2.020 0.345 2.140 1.860 ;
        RECT  1.865 0.345 2.020 0.465 ;
        RECT  1.990 1.600 2.020 1.860 ;
        RECT  1.350 1.740 1.990 1.860 ;
        RECT  1.860 0.865 1.900 1.385 ;
        RECT  1.700 1.980 1.885 2.140 ;
        RECT  1.730 0.585 1.860 1.620 ;
        RECT  1.515 0.585 1.730 0.705 ;
        RECT  1.560 1.500 1.730 1.620 ;
        RECT  0.650 1.980 1.700 2.100 ;
        RECT  1.230 0.800 1.350 1.860 ;
        RECT  0.990 0.800 1.230 0.935 ;
        RECT  0.990 1.415 1.230 1.635 ;
        RECT  0.650 1.075 1.110 1.245 ;
        RECT  0.820 0.385 0.990 0.935 ;
        RECT  0.820 1.415 0.990 1.860 ;
        RECT  0.505 0.385 0.650 2.100 ;
        RECT  0.455 0.385 0.505 0.815 ;
        RECT  0.455 1.630 0.505 2.100 ;
    END
END XNOR2X2AD
MACRO XNOR2X4AD
    CLASS CORE ;
    FOREIGN XNOR2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.270 0.510 4.410 1.810 ;
        RECT  3.265 0.510 4.270 0.640 ;
        RECT  4.000 1.640 4.270 1.810 ;
        RECT  3.875 1.640 4.000 1.920 ;
        RECT  3.385 1.800 3.875 1.920 ;
        RECT  3.265 1.800 3.385 2.135 ;
        RECT  3.095 0.380 3.265 0.810 ;
        RECT  1.505 2.015 3.265 2.135 ;
        RECT  2.515 0.690 3.095 0.810 ;
        RECT  2.300 0.620 2.515 0.810 ;
        RECT  1.765 0.620 2.300 0.740 ;
        RECT  1.595 0.620 1.765 0.790 ;
        END
        AntennaDiffArea 1.023 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.225 1.075 0.545 1.245 ;
        RECT  0.070 1.075 0.225 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.080 1.155 1.535 1.325 ;
        RECT  0.910 0.860 1.080 1.325 ;
        END
        AntennaGateArea 0.3933 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.370 -0.210 4.480 0.210 ;
        RECT  4.110 -0.210 4.370 0.390 ;
        RECT  3.650 -0.210 4.110 0.210 ;
        RECT  3.390 -0.210 3.650 0.390 ;
        RECT  1.050 -0.210 3.390 0.210 ;
        RECT  0.790 -0.210 1.050 0.390 ;
        RECT  0.265 -0.210 0.790 0.210 ;
        RECT  0.095 -0.210 0.265 0.875 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.380 2.310 4.480 2.730 ;
        RECT  4.195 1.940 4.380 2.730 ;
        RECT  3.695 2.310 4.195 2.730 ;
        RECT  3.510 2.060 3.695 2.730 ;
        RECT  1.050 2.310 3.510 2.730 ;
        RECT  0.790 2.010 1.050 2.730 ;
        RECT  0.265 2.310 0.790 2.730 ;
        RECT  0.095 1.610 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
        LAYER M1 ;
        RECT  3.965 1.400 4.060 1.520 ;
        RECT  3.965 0.760 4.010 0.880 ;
        RECT  3.740 0.760 3.965 1.520 ;
        RECT  3.700 0.760 3.740 1.050 ;
        RECT  2.905 0.930 3.700 1.050 ;
        RECT  3.250 1.185 3.420 1.625 ;
        RECT  3.145 1.455 3.250 1.625 ;
        RECT  3.025 1.455 3.145 1.890 ;
        RECT  0.790 1.770 3.025 1.890 ;
        RECT  2.680 0.380 2.940 0.570 ;
        RECT  2.785 0.930 2.905 1.635 ;
        RECT  2.180 0.930 2.785 1.050 ;
        RECT  2.645 1.515 2.785 1.635 ;
        RECT  1.365 0.380 2.680 0.500 ;
        RECT  2.495 1.175 2.665 1.380 ;
        RECT  1.800 1.260 2.495 1.380 ;
        RECT  1.920 0.860 2.180 1.050 ;
        RECT  1.680 0.910 1.800 1.650 ;
        RECT  1.460 0.910 1.680 1.030 ;
        RECT  1.170 1.530 1.680 1.650 ;
        RECT  1.340 0.760 1.460 1.030 ;
        RECT  1.245 0.380 1.365 0.630 ;
        RECT  1.200 0.760 1.340 0.880 ;
        RECT  0.790 0.510 1.245 0.630 ;
        RECT  0.670 0.510 0.790 1.890 ;
        RECT  0.635 0.510 0.670 0.875 ;
        RECT  0.635 1.610 0.670 1.890 ;
        RECT  0.465 0.445 0.635 0.875 ;
        RECT  0.465 1.610 0.635 2.040 ;
    END
END XNOR2X4AD
MACRO XNOR2XLAD
    CLASS CORE ;
    FOREIGN XNOR2XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.550 0.350 1.655 0.490 ;
        RECT  1.430 0.350 1.550 1.825 ;
        RECT  1.145 0.350 1.430 0.680 ;
        RECT  1.200 1.705 1.430 1.825 ;
        END
        AntennaDiffArea 0.11 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.380 0.865 0.770 1.105 ;
        END
        AntennaGateArea 0.0613 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.200 1.705 0.490 2.170 ;
        END
        AntennaGateArea 0.0887 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.125 -0.210 2.240 0.210 ;
        RECT  2.005 -0.210 2.125 0.420 ;
        RECT  0.635 -0.210 2.005 0.210 ;
        RECT  0.465 -0.210 0.635 0.705 ;
        RECT  0.000 -0.210 0.465 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.140 2.310 2.240 2.730 ;
        RECT  1.880 2.220 2.140 2.730 ;
        RECT  0.730 2.310 1.880 2.730 ;
        RECT  0.610 1.465 0.730 2.730 ;
        RECT  0.420 1.465 0.610 1.585 ;
        RECT  0.000 2.310 0.610 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.920 1.020 2.040 2.065 ;
        RECT  0.990 1.945 1.920 2.065 ;
        RECT  1.670 0.610 1.790 1.825 ;
        RECT  1.190 0.800 1.310 1.585 ;
        RECT  1.025 0.800 1.190 0.920 ;
        RECT  0.990 1.465 1.190 1.585 ;
        RECT  0.950 1.040 1.070 1.345 ;
        RECT  0.890 0.535 1.025 0.920 ;
        RECT  0.870 1.465 0.990 2.065 ;
        RECT  0.265 1.225 0.950 1.345 ;
        RECT  0.855 0.535 0.890 0.705 ;
        RECT  0.225 0.535 0.265 0.705 ;
        RECT  0.225 1.225 0.265 1.555 ;
        RECT  0.095 0.535 0.225 1.555 ;
    END
END XNOR2XLAD
MACRO XNOR3X1AD
    CLASS CORE ;
    FOREIGN XNOR3X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.190 0.655 5.250 1.645 ;
        RECT  5.110 0.655 5.190 1.990 ;
        RECT  5.070 0.655 5.110 0.915 ;
        RECT  5.070 1.470 5.110 1.990 ;
        END
        AntennaDiffArea 0.216 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.225 1.750 4.485 2.190 ;
        END
        AntennaGateArea 0.1345 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.865 2.750 1.405 ;
        END
        AntennaGateArea 0.1585 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.075 0.370 1.245 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.14 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.860 -0.210 5.320 0.210 ;
        RECT  4.600 -0.210 4.860 0.315 ;
        RECT  2.920 -0.210 4.600 0.210 ;
        RECT  2.730 -0.210 2.920 0.525 ;
        RECT  1.900 -0.210 2.730 0.210 ;
        RECT  1.730 -0.210 1.900 0.865 ;
        RECT  0.270 -0.210 1.730 0.210 ;
        RECT  0.100 -0.210 0.270 0.665 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.850 2.310 5.320 2.730 ;
        RECT  4.665 1.470 4.850 2.730 ;
        RECT  3.020 2.310 4.665 2.730 ;
        RECT  2.760 2.105 3.020 2.730 ;
        RECT  1.875 2.310 2.760 2.730 ;
        RECT  1.615 2.105 1.875 2.730 ;
        RECT  0.245 2.310 1.615 2.730 ;
        RECT  0.100 1.545 0.245 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.320 2.520 ;
        LAYER M1 ;
        RECT  4.865 1.000 4.930 1.260 ;
        RECT  4.745 0.455 4.865 1.260 ;
        RECT  3.685 0.455 4.745 0.575 ;
        RECT  4.350 0.735 4.415 0.905 ;
        RECT  4.350 1.375 4.415 1.545 ;
        RECT  4.230 0.735 4.350 1.545 ;
        RECT  4.200 1.005 4.230 1.545 ;
        RECT  4.045 1.005 4.200 1.265 ;
        RECT  3.925 0.695 4.110 0.815 ;
        RECT  4.020 1.725 4.090 1.985 ;
        RECT  3.925 1.385 4.020 1.985 ;
        RECT  3.900 0.695 3.925 1.985 ;
        RECT  3.805 0.695 3.900 1.505 ;
        RECT  3.090 1.865 3.900 1.985 ;
        RECT  3.685 1.625 3.780 1.745 ;
        RECT  3.515 0.455 3.685 1.745 ;
        RECT  3.210 0.410 3.330 1.680 ;
        RECT  3.150 0.410 3.210 0.670 ;
        RECT  2.970 0.960 3.090 1.985 ;
        RECT  0.860 1.865 2.970 1.985 ;
        RECT  2.470 1.625 2.640 1.745 ;
        RECT  2.470 0.355 2.535 0.525 ;
        RECT  2.350 0.355 2.470 1.745 ;
        RECT  1.100 1.625 2.350 1.745 ;
        RECT  2.110 0.640 2.230 1.505 ;
        RECT  2.060 1.335 2.110 1.505 ;
        RECT  1.340 1.385 2.060 1.505 ;
        RECT  1.610 1.025 1.930 1.195 ;
        RECT  1.490 0.380 1.610 1.195 ;
        RECT  0.610 0.380 1.490 0.500 ;
        RECT  1.340 0.645 1.370 0.905 ;
        RECT  1.220 0.645 1.340 1.505 ;
        RECT  0.980 0.990 1.100 1.745 ;
        RECT  0.860 0.620 1.060 0.740 ;
        RECT  0.740 0.620 0.860 1.985 ;
        RECT  0.490 0.380 0.610 2.045 ;
    END
END XNOR3X1AD
MACRO XNOR3X2AD
    CLASS CORE ;
    FOREIGN XNOR3X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.215 0.745 5.250 1.655 ;
        RECT  5.110 0.365 5.215 2.080 ;
        RECT  5.070 0.365 5.110 0.885 ;
        RECT  5.070 1.480 5.110 2.080 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.470 1.000 4.690 1.400 ;
        END
        AntennaGateArea 0.1826 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.900 2.750 1.420 ;
        END
        AntennaGateArea 0.1871 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.075 0.370 1.245 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.16 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.900 -0.210 5.320 0.210 ;
        RECT  4.640 -0.210 4.900 0.390 ;
        RECT  2.925 -0.210 4.640 0.210 ;
        RECT  2.755 -0.210 2.925 0.775 ;
        RECT  1.885 -0.210 2.755 0.210 ;
        RECT  1.715 -0.210 1.885 0.895 ;
        RECT  0.265 -0.210 1.715 0.210 ;
        RECT  0.095 -0.210 0.265 0.725 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.865 2.310 5.320 2.730 ;
        RECT  4.680 1.560 4.865 2.730 ;
        RECT  3.030 2.310 4.680 2.730 ;
        RECT  2.770 2.130 3.030 2.730 ;
        RECT  1.870 2.310 2.770 2.730 ;
        RECT  1.610 2.130 1.870 2.730 ;
        RECT  0.290 2.310 1.610 2.730 ;
        RECT  0.105 1.550 0.290 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.320 2.520 ;
        LAYER M1 ;
        RECT  4.830 0.510 4.950 1.265 ;
        RECT  3.650 0.510 4.830 0.630 ;
        RECT  4.350 0.760 4.520 0.880 ;
        RECT  4.350 1.565 4.445 1.735 ;
        RECT  4.230 0.760 4.350 1.735 ;
        RECT  4.035 1.070 4.230 1.210 ;
        RECT  3.935 1.350 4.105 2.010 ;
        RECT  3.915 0.760 4.100 0.880 ;
        RECT  3.915 1.350 3.935 1.470 ;
        RECT  3.090 1.890 3.935 2.010 ;
        RECT  3.795 0.760 3.915 1.470 ;
        RECT  3.650 1.600 3.735 1.770 ;
        RECT  3.530 0.510 3.650 1.770 ;
        RECT  3.210 0.345 3.330 1.770 ;
        RECT  3.125 0.345 3.210 0.775 ;
        RECT  2.970 0.960 3.090 2.010 ;
        RECT  0.860 1.890 2.970 2.010 ;
        RECT  2.470 0.605 2.565 0.775 ;
        RECT  2.470 1.560 2.565 1.730 ;
        RECT  2.350 0.605 2.470 1.770 ;
        RECT  1.100 1.650 2.350 1.770 ;
        RECT  2.100 0.635 2.230 1.530 ;
        RECT  2.075 0.635 2.100 0.895 ;
        RECT  1.350 1.410 2.100 1.530 ;
        RECT  1.595 1.065 1.945 1.235 ;
        RECT  1.475 0.380 1.595 1.235 ;
        RECT  0.610 0.380 1.475 0.500 ;
        RECT  1.230 0.660 1.350 1.530 ;
        RECT  0.980 0.990 1.100 1.770 ;
        RECT  0.860 0.670 1.050 0.790 ;
        RECT  0.740 0.670 0.860 2.010 ;
        RECT  0.490 0.380 0.610 2.045 ;
    END
END XNOR3X2AD
MACRO XNOR3X4AD
    CLASS CORE ;
    FOREIGN XNOR3X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.750 0.970 5.810 1.515 ;
        RECT  5.715 0.470 5.750 1.515 ;
        RECT  5.690 0.470 5.715 2.080 ;
        RECT  5.610 0.470 5.690 2.120 ;
        RECT  5.545 0.470 5.610 0.640 ;
        RECT  5.570 1.375 5.610 2.120 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.980 1.000 5.250 1.520 ;
        END
        AntennaGateArea 0.1864 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.805 2.730 1.375 ;
        END
        AntennaGateArea 0.187 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.075 0.370 1.245 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.16 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.075 -0.210 6.160 0.210 ;
        RECT  5.905 -0.210 6.075 0.885 ;
        RECT  5.400 -0.210 5.905 0.210 ;
        RECT  5.140 -0.210 5.400 0.390 ;
        RECT  3.575 -0.210 5.140 0.210 ;
        RECT  3.405 -0.210 3.575 0.875 ;
        RECT  2.850 -0.210 3.405 0.210 ;
        RECT  2.680 -0.210 2.850 0.570 ;
        RECT  1.885 -0.210 2.680 0.210 ;
        RECT  1.715 -0.210 1.885 0.895 ;
        RECT  0.265 -0.210 1.715 0.210 ;
        RECT  0.095 -0.210 0.265 0.720 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.070 2.310 6.160 2.730 ;
        RECT  5.900 1.600 6.070 2.730 ;
        RECT  5.365 2.310 5.900 2.730 ;
        RECT  5.180 1.665 5.365 2.730 ;
        RECT  3.675 2.310 5.180 2.730 ;
        RECT  3.415 2.130 3.675 2.730 ;
        RECT  2.875 2.310 3.415 2.730 ;
        RECT  2.615 2.130 2.875 2.730 ;
        RECT  1.870 2.310 2.615 2.730 ;
        RECT  1.610 2.130 1.870 2.730 ;
        RECT  0.290 2.310 1.610 2.730 ;
        RECT  0.105 1.550 0.290 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.370 0.760 5.490 1.265 ;
        RECT  5.295 0.760 5.370 0.880 ;
        RECT  5.175 0.510 5.295 0.880 ;
        RECT  4.250 0.510 5.175 0.630 ;
        RECT  4.860 0.760 5.020 0.880 ;
        RECT  4.860 1.650 4.975 1.820 ;
        RECT  4.740 0.760 4.860 1.820 ;
        RECT  4.730 1.090 4.740 1.820 ;
        RECT  4.665 1.090 4.730 1.350 ;
        RECT  4.515 0.775 4.620 0.945 ;
        RECT  4.515 1.535 4.610 2.055 ;
        RECT  4.490 0.775 4.515 2.055 ;
        RECT  4.395 0.775 4.490 2.010 ;
        RECT  2.970 1.890 4.395 2.010 ;
        RECT  4.200 1.555 4.275 1.725 ;
        RECT  4.200 0.510 4.250 0.680 ;
        RECT  4.080 0.510 4.200 1.725 ;
        RECT  3.700 1.475 3.960 1.770 ;
        RECT  3.745 0.350 3.865 1.175 ;
        RECT  3.625 1.055 3.745 1.175 ;
        RECT  3.625 1.475 3.700 1.595 ;
        RECT  3.385 1.055 3.625 1.595 ;
        RECT  3.280 1.055 3.385 1.175 ;
        RECT  3.225 1.475 3.385 1.595 ;
        RECT  3.160 0.395 3.280 1.175 ;
        RECT  3.105 1.475 3.225 1.735 ;
        RECT  3.045 0.395 3.160 0.825 ;
        RECT  2.970 1.010 3.040 1.270 ;
        RECT  2.850 1.010 2.970 2.010 ;
        RECT  0.860 1.890 2.850 2.010 ;
        RECT  2.435 0.395 2.490 0.565 ;
        RECT  2.435 1.500 2.490 1.670 ;
        RECT  2.315 0.395 2.435 1.770 ;
        RECT  1.100 1.650 2.315 1.770 ;
        RECT  2.075 0.635 2.195 1.530 ;
        RECT  1.350 1.410 2.075 1.530 ;
        RECT  1.595 1.065 1.945 1.235 ;
        RECT  1.475 0.380 1.595 1.235 ;
        RECT  0.610 0.380 1.475 0.500 ;
        RECT  1.230 0.660 1.350 1.530 ;
        RECT  0.980 1.000 1.100 1.770 ;
        RECT  0.860 0.670 1.050 0.790 ;
        RECT  0.740 0.670 0.860 2.010 ;
        RECT  0.490 0.380 0.610 2.045 ;
    END
END XNOR3X4AD
MACRO XNOR3XLAD
    CLASS CORE ;
    FOREIGN XNOR3XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 0.735 4.690 1.655 ;
        RECT  4.485 0.735 4.550 0.905 ;
        RECT  4.475 1.485 4.550 1.655 ;
        END
        AntennaDiffArea 0.14 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.665 1.750 3.925 2.190 ;
        END
        AntennaGateArea 0.1213 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.950 2.210 1.470 ;
        END
        AntennaGateArea 0.1421 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.075 0.310 1.245 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.1075 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.330 -0.210 4.760 0.210 ;
        RECT  4.070 -0.210 4.330 0.375 ;
        RECT  2.465 -0.210 4.070 0.210 ;
        RECT  2.295 -0.210 2.465 0.415 ;
        RECT  1.905 -0.210 2.295 0.210 ;
        RECT  1.750 -0.210 1.905 0.560 ;
        RECT  0.270 -0.210 1.750 0.210 ;
        RECT  0.100 -0.210 0.270 0.740 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.310 2.310 4.760 2.730 ;
        RECT  4.095 1.455 4.310 2.730 ;
        RECT  2.520 2.310 4.095 2.730 ;
        RECT  2.260 2.150 2.520 2.730 ;
        RECT  1.880 2.310 2.260 2.730 ;
        RECT  1.620 2.105 1.880 2.730 ;
        RECT  0.255 2.310 1.620 2.730 ;
        RECT  0.085 1.625 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.760 2.520 ;
        LAYER M1 ;
        RECT  4.290 1.055 4.405 1.225 ;
        RECT  4.170 0.495 4.290 1.225 ;
        RECT  3.830 0.495 4.170 0.615 ;
        RECT  3.835 1.480 3.940 1.600 ;
        RECT  3.835 0.735 3.895 0.905 ;
        RECT  3.680 0.735 3.835 1.600 ;
        RECT  3.710 0.395 3.830 0.615 ;
        RECT  3.175 0.395 3.710 0.515 ;
        RECT  3.560 1.095 3.680 1.295 ;
        RECT  3.435 0.700 3.560 0.960 ;
        RECT  3.435 1.725 3.540 2.030 ;
        RECT  3.315 0.700 3.435 2.030 ;
        RECT  2.500 1.900 3.315 2.030 ;
        RECT  3.055 0.395 3.175 1.760 ;
        RECT  2.995 0.685 3.055 0.855 ;
        RECT  3.005 1.590 3.055 1.760 ;
        RECT  2.690 0.685 2.810 1.750 ;
        RECT  2.615 0.685 2.690 0.855 ;
        RECT  2.625 1.580 2.690 1.750 ;
        RECT  2.500 0.990 2.570 1.250 ;
        RECT  2.380 0.990 2.500 2.030 ;
        RECT  0.860 1.865 2.380 1.985 ;
        RECT  1.885 1.625 2.130 1.745 ;
        RECT  1.885 0.710 2.120 0.830 ;
        RECT  1.755 0.710 1.885 1.745 ;
        RECT  1.100 1.625 1.755 1.745 ;
        RECT  1.500 0.380 1.630 1.210 ;
        RECT  0.610 0.380 1.500 0.500 ;
        RECT  1.460 1.040 1.500 1.210 ;
        RECT  1.340 1.385 1.480 1.505 ;
        RECT  1.340 0.645 1.380 0.905 ;
        RECT  1.220 0.645 1.340 1.505 ;
        RECT  0.980 0.990 1.100 1.745 ;
        RECT  0.860 0.640 1.060 0.790 ;
        RECT  0.740 0.640 0.860 1.985 ;
        RECT  0.475 0.380 0.610 2.100 ;
    END
END XNOR3XLAD
MACRO XOR2X1AD
    CLASS CORE ;
    FOREIGN XOR2X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.530 0.350 1.655 0.490 ;
        RECT  1.410 0.350 1.530 1.825 ;
        RECT  1.145 0.350 1.410 0.670 ;
        RECT  1.160 1.705 1.410 1.825 ;
        END
        AntennaDiffArea 0.158 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 0.865 0.780 1.095 ;
        END
        AntennaGateArea 0.09 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.170 1.705 0.490 2.160 ;
        END
        AntennaGateArea 0.1073 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.130 -0.210 2.240 0.210 ;
        RECT  2.010 -0.210 2.130 0.430 ;
        RECT  0.625 -0.210 2.010 0.210 ;
        RECT  0.455 -0.210 0.625 0.700 ;
        RECT  0.000 -0.210 0.455 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.310 2.240 2.730 ;
        RECT  1.885 2.220 2.145 2.730 ;
        RECT  0.740 2.310 1.885 2.730 ;
        RECT  0.610 1.465 0.740 2.730 ;
        RECT  0.410 1.465 0.610 1.585 ;
        RECT  0.000 2.310 0.610 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.900 1.015 2.020 2.090 ;
        RECT  0.980 1.970 1.900 2.090 ;
        RECT  1.650 0.660 1.770 1.850 ;
        RECT  1.170 0.820 1.290 1.585 ;
        RECT  1.025 0.820 1.170 0.940 ;
        RECT  0.980 1.465 1.170 1.585 ;
        RECT  0.930 1.060 1.050 1.345 ;
        RECT  0.905 0.555 1.025 0.940 ;
        RECT  0.860 1.465 0.980 2.090 ;
        RECT  0.265 1.225 0.930 1.345 ;
        RECT  0.815 0.555 0.905 0.725 ;
        RECT  0.230 0.525 0.265 0.695 ;
        RECT  0.230 1.225 0.265 1.565 ;
        RECT  0.095 0.525 0.230 1.565 ;
    END
END XOR2X1AD
MACRO XOR2X2AD
    CLASS CORE ;
    FOREIGN XOR2X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 0.690 1.970 2.090 ;
        END
        AntennaDiffArea 0.506 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.065 2.730 1.375 ;
        RECT  2.450 1.065 2.590 1.240 ;
        END
        AntennaGateArea 0.162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.630 1.055 0.905 1.485 ;
        END
        AntennaGateArea 0.1902 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.715 -0.210 2.800 0.210 ;
        RECT  2.545 -0.210 2.715 0.815 ;
        RECT  0.615 -0.210 2.545 0.210 ;
        RECT  0.445 -0.210 0.615 0.675 ;
        RECT  0.000 -0.210 0.445 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.715 2.310 2.800 2.730 ;
        RECT  2.545 1.660 2.715 2.730 ;
        RECT  0.660 2.310 2.545 2.730 ;
        RECT  0.400 2.130 0.660 2.730 ;
        RECT  0.000 2.310 0.400 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.800 2.520 ;
        LAYER M1 ;
        RECT  2.330 1.660 2.355 2.090 ;
        RECT  2.210 0.420 2.330 2.090 ;
        RECT  0.855 0.420 2.210 0.540 ;
        RECT  2.185 1.660 2.210 2.090 ;
        RECT  1.395 0.690 1.515 2.090 ;
        RECT  1.345 1.660 1.395 2.090 ;
        RECT  0.230 1.890 1.345 2.010 ;
        RECT  1.200 0.970 1.250 1.230 ;
        RECT  1.080 0.660 1.200 1.770 ;
        RECT  0.975 0.660 1.080 0.920 ;
        RECT  0.810 1.650 1.080 1.770 ;
        RECT  0.735 0.420 0.855 0.920 ;
        RECT  0.470 0.800 0.735 0.920 ;
        RECT  0.350 0.800 0.470 1.300 ;
        RECT  0.110 0.395 0.230 2.010 ;
    END
END XOR2X2AD
MACRO XOR2X3AD
    CLASS CORE ;
    FOREIGN XOR2X3AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.605 1.920 3.410 2.040 ;
        RECT  3.140 0.760 3.400 0.960 ;
        RECT  2.605 0.840 3.140 0.960 ;
        RECT  2.435 0.620 2.605 0.960 ;
        RECT  2.435 1.555 2.605 2.040 ;
        RECT  1.890 0.620 2.435 0.740 ;
        RECT  1.890 1.555 2.435 1.675 ;
        RECT  1.750 0.620 1.890 1.850 ;
        RECT  1.700 0.620 1.750 0.910 ;
        RECT  1.705 1.680 1.750 1.850 ;
        END
        AntennaDiffArea 0.728 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.065 0.540 1.235 ;
        RECT  0.070 1.065 0.210 1.655 ;
        END
        AntennaGateArea 0.2444 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 0.965 1.300 1.375 ;
        END
        AntennaGateArea 0.2963 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.365 -0.210 4.480 0.210 ;
        RECT  4.180 -0.210 4.365 0.950 ;
        RECT  3.660 -0.210 4.180 0.210 ;
        RECT  3.400 -0.210 3.660 0.300 ;
        RECT  1.080 -0.210 3.400 0.210 ;
        RECT  0.820 -0.210 1.080 0.300 ;
        RECT  0.265 -0.210 0.820 0.210 ;
        RECT  0.095 -0.210 0.265 0.855 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.380 2.310 4.480 2.730 ;
        RECT  4.210 1.470 4.380 2.730 ;
        RECT  3.670 2.310 4.210 2.730 ;
        RECT  3.550 1.575 3.670 2.730 ;
        RECT  3.410 1.575 3.550 1.695 ;
        RECT  1.025 2.310 3.550 2.730 ;
        RECT  0.855 2.095 1.025 2.730 ;
        RECT  0.265 2.310 0.855 2.730 ;
        RECT  0.095 1.785 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
        LAYER M1 ;
        RECT  3.835 0.475 4.005 1.925 ;
        RECT  3.030 1.335 3.835 1.455 ;
        RECT  3.640 1.045 3.695 1.215 ;
        RECT  3.520 0.520 3.640 1.215 ;
        RECT  3.030 0.520 3.520 0.640 ;
        RECT  2.890 0.520 3.030 0.680 ;
        RECT  2.770 1.170 3.030 1.660 ;
        RECT  2.770 0.380 2.890 0.680 ;
        RECT  1.410 0.380 2.770 0.500 ;
        RECT  2.280 1.170 2.770 1.290 ;
        RECT  2.160 0.860 2.280 1.290 ;
        RECT  2.020 1.850 2.280 2.140 ;
        RECT  2.020 0.860 2.160 0.980 ;
        RECT  1.300 2.020 2.020 2.140 ;
        RECT  1.565 1.255 1.625 1.515 ;
        RECT  1.445 0.720 1.565 1.720 ;
        RECT  1.425 0.720 1.445 0.840 ;
        RECT  1.255 1.550 1.445 1.720 ;
        RECT  1.255 0.670 1.425 0.840 ;
        RECT  1.290 0.380 1.410 0.545 ;
        RECT  1.180 1.840 1.300 2.140 ;
        RECT  0.780 0.425 1.290 0.545 ;
        RECT  0.780 1.840 1.180 1.960 ;
        RECT  0.660 0.425 0.780 1.960 ;
        RECT  0.465 0.425 0.660 0.855 ;
        RECT  0.465 1.530 0.660 1.960 ;
    END
END XOR2X3AD
MACRO XOR2X4AD
    CLASS CORE ;
    FOREIGN XOR2X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.435 0.760 3.200 0.880 ;
        RECT  2.985 1.695 3.155 2.125 ;
        RECT  2.435 1.780 2.985 1.900 ;
        RECT  2.265 0.625 2.435 0.880 ;
        RECT  2.265 1.695 2.435 2.125 ;
        RECT  1.785 0.625 2.265 0.745 ;
        RECT  1.890 1.780 2.265 1.900 ;
        RECT  1.785 1.285 1.890 1.900 ;
        RECT  1.665 0.625 1.785 1.900 ;
        RECT  1.570 0.625 1.665 0.885 ;
        RECT  1.545 1.730 1.665 1.900 ;
        END
        AntennaDiffArea 1 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.075 0.545 1.245 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.324 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.065 1.125 1.235 ;
        RECT  0.910 1.065 1.050 1.675 ;
        END
        AntennaGateArea 0.3893 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.285 -0.210 4.480 0.210 ;
        RECT  4.115 -0.210 4.285 0.800 ;
        RECT  3.590 -0.210 4.115 0.210 ;
        RECT  3.330 -0.210 3.590 0.390 ;
        RECT  1.030 -0.210 3.330 0.210 ;
        RECT  0.770 -0.210 1.030 0.390 ;
        RECT  0.265 -0.210 0.770 0.210 ;
        RECT  0.095 -0.210 0.265 0.715 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.285 2.310 4.480 2.730 ;
        RECT  4.115 1.690 4.285 2.730 ;
        RECT  3.545 2.310 4.115 2.730 ;
        RECT  3.375 1.690 3.545 2.730 ;
        RECT  0.985 2.310 3.375 2.730 ;
        RECT  0.815 2.105 0.985 2.730 ;
        RECT  0.265 2.310 0.815 2.730 ;
        RECT  0.095 1.555 0.265 2.730 ;
        RECT  0.000 2.310 0.095 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.480 2.520 ;
        LAYER M1 ;
        RECT  3.745 0.370 3.915 2.125 ;
        RECT  2.840 1.430 3.745 1.550 ;
        RECT  3.535 1.050 3.585 1.220 ;
        RECT  3.415 0.520 3.535 1.220 ;
        RECT  2.840 0.520 3.415 0.640 ;
        RECT  2.580 0.380 2.840 0.640 ;
        RECT  2.735 1.430 2.840 1.650 ;
        RECT  2.580 1.080 2.735 1.650 ;
        RECT  1.290 0.380 2.580 0.500 ;
        RECT  2.130 1.080 2.580 1.200 ;
        RECT  1.990 0.865 2.130 1.200 ;
        RECT  1.245 2.020 2.120 2.140 ;
        RECT  1.905 0.865 1.990 1.035 ;
        RECT  1.410 1.135 1.500 1.305 ;
        RECT  1.290 0.760 1.410 1.675 ;
        RECT  1.170 0.380 1.290 0.630 ;
        RECT  1.150 0.760 1.290 0.880 ;
        RECT  1.195 1.505 1.290 1.675 ;
        RECT  1.125 1.865 1.245 2.140 ;
        RECT  0.785 0.510 1.170 0.630 ;
        RECT  0.785 1.865 1.125 1.985 ;
        RECT  0.665 0.510 0.785 1.985 ;
        RECT  0.625 0.510 0.665 0.835 ;
        RECT  0.455 1.555 0.665 1.985 ;
        RECT  0.455 0.405 0.625 0.835 ;
    END
END XOR2X4AD
MACRO XOR2X8AD
    CLASS CORE ;
    FOREIGN XOR2X8AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.505 0.760 5.990 0.880 ;
        RECT  5.775 1.695 5.945 2.130 ;
        RECT  5.225 1.790 5.775 2.130 ;
        RECT  5.055 1.695 5.225 2.130 ;
        RECT  4.505 1.790 5.055 2.130 ;
        RECT  4.335 0.625 4.505 0.880 ;
        RECT  4.335 1.520 4.505 2.130 ;
        RECT  3.090 0.625 4.335 0.770 ;
        RECT  3.710 1.520 4.335 1.850 ;
        RECT  3.290 1.280 3.710 1.850 ;
        RECT  3.090 1.280 3.290 1.680 ;
        RECT  2.895 0.625 3.090 1.680 ;
        END
        AntennaDiffArea 1.708 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.825 1.075 1.340 1.375 ;
        END
        AntennaGateArea 0.648 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.415 0.810 2.740 1.095 ;
        RECT  2.240 0.810 2.415 1.245 ;
        RECT  2.025 1.075 2.240 1.245 ;
        END
        AntennaGateArea 0.7777 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.745 -0.210 7.840 0.210 ;
        RECT  7.575 -0.210 7.745 0.800 ;
        RECT  7.005 -0.210 7.575 0.210 ;
        RECT  6.835 -0.210 7.005 0.800 ;
        RECT  6.330 -0.210 6.835 0.210 ;
        RECT  6.070 -0.210 6.330 0.390 ;
        RECT  2.500 -0.210 6.070 0.210 ;
        RECT  2.240 -0.210 2.500 0.390 ;
        RECT  1.740 -0.210 2.240 0.210 ;
        RECT  1.480 -0.210 1.740 0.390 ;
        RECT  0.975 -0.210 1.480 0.210 ;
        RECT  0.805 -0.210 0.975 0.435 ;
        RECT  0.255 -0.210 0.805 0.210 ;
        RECT  0.085 -0.210 0.255 0.715 ;
        RECT  0.000 -0.210 0.085 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  7.745 2.310 7.840 2.730 ;
        RECT  7.575 1.690 7.745 2.730 ;
        RECT  7.005 2.310 7.575 2.730 ;
        RECT  6.835 1.690 7.005 2.730 ;
        RECT  6.285 2.310 6.835 2.730 ;
        RECT  6.115 1.690 6.285 2.730 ;
        RECT  2.455 2.310 6.115 2.730 ;
        RECT  2.285 2.105 2.455 2.730 ;
        RECT  1.695 2.310 2.285 2.730 ;
        RECT  1.525 2.105 1.695 2.730 ;
        RECT  0.975 2.310 1.525 2.730 ;
        RECT  0.805 1.845 0.975 2.730 ;
        RECT  0.255 2.310 0.805 2.730 ;
        RECT  0.085 1.460 0.255 2.730 ;
        RECT  0.000 2.310 0.085 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 7.840 2.520 ;
        LAYER M1 ;
        RECT  7.205 0.370 7.375 2.125 ;
        RECT  6.645 1.365 7.205 1.550 ;
        RECT  6.475 0.370 6.645 2.125 ;
        RECT  5.630 1.365 6.475 1.550 ;
        RECT  6.230 1.050 6.355 1.220 ;
        RECT  6.110 0.520 6.230 1.220 ;
        RECT  4.910 0.520 6.110 0.640 ;
        RECT  5.925 1.050 6.110 1.220 ;
        RECT  5.370 1.365 5.630 1.650 ;
        RECT  4.910 1.365 5.370 1.550 ;
        RECT  4.650 0.380 4.910 0.640 ;
        RECT  4.650 1.080 4.910 1.650 ;
        RECT  2.740 0.380 4.650 0.500 ;
        RECT  4.200 1.080 4.650 1.250 ;
        RECT  4.060 0.890 4.200 1.250 ;
        RECT  3.040 2.020 4.190 2.140 ;
        RECT  3.210 0.890 4.060 1.035 ;
        RECT  2.920 1.815 3.040 2.140 ;
        RECT  1.600 1.815 2.920 1.985 ;
        RECT  2.585 1.215 2.755 1.645 ;
        RECT  2.620 0.380 2.740 0.630 ;
        RECT  1.600 0.510 2.620 0.630 ;
        RECT  2.075 1.385 2.585 1.505 ;
        RECT  1.905 0.760 2.120 0.880 ;
        RECT  1.905 1.385 2.075 1.675 ;
        RECT  1.785 0.760 1.905 1.675 ;
        RECT  1.480 0.510 1.600 1.985 ;
        RECT  1.335 0.510 1.480 0.835 ;
        RECT  1.335 1.590 1.480 1.985 ;
        RECT  1.165 0.405 1.335 0.835 ;
        RECT  1.165 1.590 1.335 2.020 ;
        RECT  0.615 0.605 1.165 0.725 ;
        RECT  0.615 1.590 1.165 1.710 ;
        RECT  0.590 0.405 0.615 0.835 ;
        RECT  0.590 1.460 0.615 2.150 ;
        RECT  0.470 0.405 0.590 2.150 ;
        RECT  0.445 0.405 0.470 0.835 ;
        RECT  0.445 1.460 0.470 2.150 ;
    END
END XOR2X8AD
MACRO XOR2XLAD
    CLASS CORE ;
    FOREIGN XOR2XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.530 0.350 1.655 0.490 ;
        RECT  1.410 0.350 1.530 1.825 ;
        RECT  1.145 0.350 1.410 0.665 ;
        RECT  1.200 1.705 1.410 1.825 ;
        END
        AntennaDiffArea 0.138 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.865 0.780 1.095 ;
        END
        AntennaGateArea 0.06 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.705 0.490 2.150 ;
        RECT  0.110 1.890 0.350 2.150 ;
        END
        AntennaGateArea 0.0894 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.130 -0.210 2.240 0.210 ;
        RECT  2.010 -0.210 2.130 0.425 ;
        RECT  0.625 -0.210 2.010 0.210 ;
        RECT  0.455 -0.210 0.625 0.690 ;
        RECT  0.000 -0.210 0.455 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  2.170 2.310 2.240 2.730 ;
        RECT  1.910 2.220 2.170 2.730 ;
        RECT  0.740 2.310 1.910 2.730 ;
        RECT  0.610 1.465 0.740 2.730 ;
        RECT  0.410 1.465 0.610 1.585 ;
        RECT  0.000 2.310 0.610 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 2.240 2.520 ;
        LAYER M1 ;
        RECT  1.900 1.015 2.020 2.100 ;
        RECT  0.980 1.980 1.900 2.100 ;
        RECT  1.660 0.610 1.780 1.860 ;
        RECT  1.170 0.785 1.290 1.585 ;
        RECT  1.025 0.785 1.170 0.905 ;
        RECT  0.980 1.465 1.170 1.585 ;
        RECT  0.930 1.025 1.050 1.345 ;
        RECT  0.905 0.520 1.025 0.905 ;
        RECT  0.860 1.465 0.980 2.100 ;
        RECT  0.265 1.225 0.930 1.345 ;
        RECT  0.815 0.520 0.905 0.690 ;
        RECT  0.230 0.520 0.265 0.690 ;
        RECT  0.230 1.225 0.265 1.545 ;
        RECT  0.095 0.520 0.230 1.545 ;
    END
END XOR2XLAD
MACRO XOR3X1AD
    CLASS CORE ;
    FOREIGN XOR3X1AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.110 0.685 5.250 1.990 ;
        RECT  5.065 0.685 5.110 0.855 ;
        RECT  5.080 1.470 5.110 1.990 ;
        END
        AntennaDiffArea 0.216 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.225 1.750 4.455 2.185 ;
        END
        AntennaGateArea 0.1284 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.865 2.745 1.495 ;
        END
        AntennaGateArea 0.1582 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.075 0.370 1.245 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.14 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.860 -0.210 5.320 0.210 ;
        RECT  4.600 -0.210 4.860 0.315 ;
        RECT  2.920 -0.210 4.600 0.210 ;
        RECT  2.735 -0.210 2.920 0.530 ;
        RECT  1.890 -0.210 2.735 0.210 ;
        RECT  1.720 -0.210 1.890 0.870 ;
        RECT  0.265 -0.210 1.720 0.210 ;
        RECT  0.095 -0.210 0.265 0.665 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.850 2.310 5.320 2.730 ;
        RECT  4.665 1.470 4.850 2.730 ;
        RECT  3.010 2.310 4.665 2.730 ;
        RECT  2.750 2.210 3.010 2.730 ;
        RECT  1.870 2.310 2.750 2.730 ;
        RECT  1.610 2.105 1.870 2.730 ;
        RECT  0.245 2.310 1.610 2.730 ;
        RECT  0.100 1.550 0.245 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.320 2.520 ;
        LAYER M1 ;
        RECT  4.865 1.005 4.930 1.265 ;
        RECT  4.745 0.455 4.865 1.265 ;
        RECT  4.390 0.455 4.745 0.575 ;
        RECT  4.285 0.735 4.455 1.590 ;
        RECT  4.240 0.380 4.390 0.575 ;
        RECT  4.035 0.985 4.285 1.245 ;
        RECT  3.675 0.380 4.240 0.500 ;
        RECT  3.915 0.625 4.120 0.745 ;
        RECT  4.035 1.675 4.105 2.020 ;
        RECT  3.915 1.385 4.035 2.020 ;
        RECT  3.795 0.625 3.915 1.505 ;
        RECT  3.065 1.880 3.915 2.020 ;
        RECT  3.675 1.625 3.795 1.745 ;
        RECT  3.505 0.380 3.675 1.745 ;
        RECT  3.235 0.455 3.355 1.760 ;
        RECT  3.125 0.455 3.235 0.625 ;
        RECT  3.185 1.590 3.235 1.760 ;
        RECT  3.065 0.900 3.110 1.420 ;
        RECT  2.945 0.900 3.065 2.020 ;
        RECT  0.860 1.865 2.945 1.985 ;
        RECT  2.470 1.625 2.615 1.745 ;
        RECT  2.470 0.385 2.580 0.505 ;
        RECT  2.350 0.385 2.470 1.745 ;
        RECT  2.320 0.385 2.350 0.505 ;
        RECT  1.100 1.625 2.350 1.745 ;
        RECT  2.060 0.640 2.230 1.505 ;
        RECT  1.360 1.385 2.060 1.505 ;
        RECT  1.600 1.015 1.685 1.185 ;
        RECT  1.480 0.400 1.600 1.185 ;
        RECT  0.610 0.400 1.480 0.520 ;
        RECT  1.220 0.645 1.360 1.505 ;
        RECT  0.980 0.990 1.100 1.745 ;
        RECT  0.860 0.640 1.060 0.760 ;
        RECT  0.740 0.640 0.860 1.985 ;
        RECT  0.490 0.400 0.610 2.045 ;
    END
END XOR3X1AD
MACRO XOR3X2AD
    CLASS CORE ;
    FOREIGN XOR3X2AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.110 0.360 5.250 2.000 ;
        RECT  5.080 0.360 5.110 0.880 ;
        RECT  5.080 1.480 5.110 2.000 ;
        END
        AntennaDiffArea 0.373 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.240 1.705 4.500 2.185 ;
        END
        AntennaGateArea 0.1841 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.590 0.995 2.760 1.445 ;
        END
        AntennaGateArea 0.1874 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.075 0.350 1.245 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.16 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.890 -0.210 5.320 0.210 ;
        RECT  4.730 -0.210 4.890 0.810 ;
        RECT  2.945 -0.210 4.730 0.210 ;
        RECT  2.775 -0.210 2.945 0.795 ;
        RECT  1.875 -0.210 2.775 0.210 ;
        RECT  1.705 -0.210 1.875 0.865 ;
        RECT  0.270 -0.210 1.705 0.210 ;
        RECT  0.100 -0.210 0.270 0.665 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.885 2.310 5.320 2.730 ;
        RECT  4.690 1.480 4.885 2.730 ;
        RECT  3.010 2.310 4.690 2.730 ;
        RECT  2.750 2.210 3.010 2.730 ;
        RECT  1.875 2.310 2.750 2.730 ;
        RECT  1.615 2.130 1.875 2.730 ;
        RECT  0.245 2.310 1.615 2.730 ;
        RECT  0.100 1.550 0.245 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 5.320 2.520 ;
        LAYER M1 ;
        RECT  4.610 0.990 4.990 1.250 ;
        RECT  4.490 0.395 4.610 1.250 ;
        RECT  3.665 0.395 4.490 0.515 ;
        RECT  4.370 1.375 4.455 1.545 ;
        RECT  4.220 0.635 4.370 1.545 ;
        RECT  4.210 0.970 4.220 1.545 ;
        RECT  4.035 0.970 4.210 1.230 ;
        RECT  3.915 0.650 4.090 0.770 ;
        RECT  3.940 1.365 4.060 2.010 ;
        RECT  3.915 1.365 3.940 1.485 ;
        RECT  3.065 1.865 3.940 2.010 ;
        RECT  3.795 0.650 3.915 1.485 ;
        RECT  3.665 1.625 3.770 1.745 ;
        RECT  3.495 0.365 3.665 1.745 ;
        RECT  3.235 0.365 3.355 1.730 ;
        RECT  3.135 0.365 3.235 0.795 ;
        RECT  3.185 1.560 3.235 1.730 ;
        RECT  3.065 0.945 3.090 1.205 ;
        RECT  2.970 0.945 3.065 2.010 ;
        RECT  2.945 0.985 2.970 2.010 ;
        RECT  0.830 1.890 2.945 2.010 ;
        RECT  2.470 1.600 2.580 1.770 ;
        RECT  2.470 0.685 2.550 0.855 ;
        RECT  2.350 0.625 2.470 1.770 ;
        RECT  1.070 1.650 2.350 1.770 ;
        RECT  2.180 1.410 2.230 1.530 ;
        RECT  2.180 0.650 2.210 0.820 ;
        RECT  2.010 0.650 2.180 1.530 ;
        RECT  1.335 1.410 2.010 1.530 ;
        RECT  1.585 1.065 1.685 1.235 ;
        RECT  1.465 0.380 1.585 1.235 ;
        RECT  0.590 0.380 1.465 0.500 ;
        RECT  1.190 0.645 1.335 1.530 ;
        RECT  1.165 0.645 1.190 0.815 ;
        RECT  0.950 1.000 1.070 1.770 ;
        RECT  0.830 0.670 1.020 0.825 ;
        RECT  0.760 0.670 0.830 2.010 ;
        RECT  0.710 0.705 0.760 2.010 ;
        RECT  0.470 0.340 0.590 2.045 ;
    END
END XOR3X2AD
MACRO XOR3X4AD
    CLASS CORE ;
    FOREIGN XOR3X4AD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.750 0.970 5.810 1.515 ;
        RECT  5.715 0.350 5.750 1.515 ;
        RECT  5.610 0.350 5.715 2.075 ;
        RECT  5.545 0.350 5.610 0.780 ;
        RECT  5.545 1.380 5.610 2.075 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.100 1.145 5.250 1.520 ;
        RECT  4.980 1.000 5.100 1.520 ;
        END
        AntennaGateArea 0.1874 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.555 0.805 2.730 1.375 ;
        END
        AntennaGateArea 0.187 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.075 0.370 1.245 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.16 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.075 -0.210 6.160 0.210 ;
        RECT  5.905 -0.210 6.075 0.885 ;
        RECT  5.400 -0.210 5.905 0.210 ;
        RECT  5.140 -0.210 5.400 0.390 ;
        RECT  3.575 -0.210 5.140 0.210 ;
        RECT  3.405 -0.210 3.575 0.875 ;
        RECT  2.850 -0.210 3.405 0.210 ;
        RECT  2.680 -0.210 2.850 0.570 ;
        RECT  1.870 -0.210 2.680 0.210 ;
        RECT  1.700 -0.210 1.870 0.895 ;
        RECT  0.265 -0.210 1.700 0.210 ;
        RECT  0.095 -0.210 0.265 0.720 ;
        RECT  0.000 -0.210 0.095 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  6.070 2.310 6.160 2.730 ;
        RECT  5.900 1.600 6.070 2.730 ;
        RECT  5.365 2.310 5.900 2.730 ;
        RECT  5.180 1.665 5.365 2.730 ;
        RECT  3.675 2.310 5.180 2.730 ;
        RECT  3.415 2.130 3.675 2.730 ;
        RECT  2.875 2.310 3.415 2.730 ;
        RECT  2.615 2.130 2.875 2.730 ;
        RECT  1.870 2.310 2.615 2.730 ;
        RECT  1.610 2.130 1.870 2.730 ;
        RECT  0.290 2.310 1.610 2.730 ;
        RECT  0.105 1.550 0.290 2.730 ;
        RECT  0.000 2.310 0.105 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 6.160 2.520 ;
        LAYER M1 ;
        RECT  5.395 0.905 5.490 1.265 ;
        RECT  5.370 0.510 5.395 1.265 ;
        RECT  5.275 0.510 5.370 1.025 ;
        RECT  4.995 0.510 5.275 0.630 ;
        RECT  4.860 0.760 5.090 0.880 ;
        RECT  4.875 0.385 4.995 0.630 ;
        RECT  4.860 1.650 4.975 1.820 ;
        RECT  4.260 0.385 4.875 0.505 ;
        RECT  4.740 0.760 4.860 1.820 ;
        RECT  4.665 0.970 4.740 1.230 ;
        RECT  4.515 0.625 4.620 0.795 ;
        RECT  4.515 1.440 4.620 2.010 ;
        RECT  4.395 0.625 4.515 2.010 ;
        RECT  2.970 1.890 4.395 2.010 ;
        RECT  4.140 0.385 4.260 1.725 ;
        RECT  4.060 0.510 4.140 0.680 ;
        RECT  4.090 1.555 4.140 1.725 ;
        RECT  3.685 1.475 3.945 1.770 ;
        RECT  3.725 0.350 3.845 1.175 ;
        RECT  3.625 1.055 3.725 1.175 ;
        RECT  3.625 1.475 3.685 1.595 ;
        RECT  3.385 1.055 3.625 1.595 ;
        RECT  3.280 1.055 3.385 1.175 ;
        RECT  3.225 1.475 3.385 1.595 ;
        RECT  3.160 0.395 3.280 1.175 ;
        RECT  3.105 1.475 3.225 1.735 ;
        RECT  3.045 0.395 3.160 0.825 ;
        RECT  2.970 1.010 3.040 1.270 ;
        RECT  2.850 1.010 2.970 2.010 ;
        RECT  0.860 1.890 2.850 2.010 ;
        RECT  2.425 0.395 2.480 0.565 ;
        RECT  2.425 1.500 2.480 1.670 ;
        RECT  2.305 0.395 2.425 1.770 ;
        RECT  1.100 1.650 2.305 1.770 ;
        RECT  2.060 0.690 2.185 1.530 ;
        RECT  1.340 1.410 2.060 1.530 ;
        RECT  1.580 1.020 1.920 1.280 ;
        RECT  1.460 0.380 1.580 1.280 ;
        RECT  0.610 0.380 1.460 0.500 ;
        RECT  1.220 0.660 1.340 1.530 ;
        RECT  0.980 1.000 1.100 1.770 ;
        RECT  0.860 0.670 1.050 0.790 ;
        RECT  0.740 0.670 0.860 2.010 ;
        RECT  0.490 0.340 0.610 2.045 ;
    END
END XOR3X4AD
MACRO XOR3XLAD
    CLASS CORE ;
    FOREIGN XOR3XLAD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.760 BY 2.520 ;
    SYMMETRY X Y ;
    SITE TSM90NMADSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 0.695 4.690 1.670 ;
        RECT  4.495 0.695 4.550 0.865 ;
        RECT  4.520 1.410 4.550 1.670 ;
        END
        AntennaDiffArea 0.148 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.665 1.750 3.945 2.190 ;
        END
        AntennaGateArea 0.1148 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.030 0.920 2.225 1.375 ;
        END
        AntennaGateArea 0.1431 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.210 1.030 0.330 1.290 ;
        RECT  0.070 0.865 0.210 1.375 ;
        END
        AntennaGateArea 0.1075 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.340 -0.210 4.760 0.210 ;
        RECT  4.080 -0.210 4.340 0.315 ;
        RECT  2.495 -0.210 4.080 0.210 ;
        RECT  2.325 -0.210 2.495 0.370 ;
        RECT  1.895 -0.210 2.325 0.210 ;
        RECT  1.740 -0.210 1.895 0.485 ;
        RECT  0.270 -0.210 1.740 0.210 ;
        RECT  0.100 -0.210 0.270 0.720 ;
        RECT  0.000 -0.210 0.100 0.210 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  4.330 2.310 4.760 2.730 ;
        RECT  4.125 1.380 4.330 2.730 ;
        RECT  4.070 1.380 4.125 1.580 ;
        RECT  2.540 2.310 4.125 2.730 ;
        RECT  2.280 2.120 2.540 2.730 ;
        RECT  1.870 2.310 2.280 2.730 ;
        RECT  1.610 2.120 1.870 2.730 ;
        RECT  0.245 2.310 1.610 2.730 ;
        RECT  0.100 1.550 0.245 2.730 ;
        RECT  0.000 2.310 0.100 2.730 ;
        END
    END VDD
	 OBS
	 LAYER RVT ;
	 RECT 0 0 4.760 2.520 ;
        LAYER M1 ;
        RECT  4.320 0.995 4.390 1.255 ;
        RECT  4.200 0.455 4.320 1.255 ;
        RECT  3.830 0.455 4.200 0.575 ;
        RECT  3.865 1.385 3.915 1.555 ;
        RECT  3.865 0.695 3.905 0.865 ;
        RECT  3.715 0.695 3.865 1.555 ;
        RECT  3.710 0.380 3.830 0.575 ;
        RECT  3.560 1.000 3.715 1.190 ;
        RECT  3.185 0.380 3.710 0.500 ;
        RECT  3.435 0.620 3.545 0.790 ;
        RECT  3.435 1.340 3.540 1.860 ;
        RECT  3.315 0.620 3.435 2.000 ;
        RECT  2.500 1.880 3.315 2.000 ;
        RECT  3.015 0.380 3.185 1.730 ;
        RECT  2.720 0.630 2.840 1.720 ;
        RECT  2.645 0.630 2.720 0.800 ;
        RECT  2.645 1.550 2.720 1.720 ;
        RECT  2.500 0.980 2.580 1.240 ;
        RECT  2.380 0.980 2.500 2.000 ;
        RECT  0.860 1.880 2.380 2.000 ;
        RECT  1.885 1.510 2.160 1.715 ;
        RECT  1.885 0.630 2.105 0.800 ;
        RECT  1.755 0.630 1.885 1.760 ;
        RECT  1.100 1.640 1.755 1.760 ;
        RECT  1.500 0.380 1.620 1.255 ;
        RECT  0.610 0.380 1.500 0.500 ;
        RECT  1.340 1.400 1.480 1.520 ;
        RECT  1.340 0.645 1.380 0.905 ;
        RECT  1.220 0.645 1.340 1.520 ;
        RECT  0.980 0.990 1.100 1.760 ;
        RECT  0.860 0.650 1.060 0.770 ;
        RECT  0.740 0.650 0.860 2.000 ;
        RECT  0.475 0.380 0.610 2.070 ;
    END
END XOR3XLAD

END LIBRARY
